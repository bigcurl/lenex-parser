<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0"><CONSTRUCTOR name="MSECM(R) Export Module" registration="Turnerbund 1888 Erlangen e.V. Schwimmabteilung" version="6.2023.117"><CONTACT city="Hoehenkirchen" country="GER" email="info@msecm.com" fax="+49 8102 748084" internet="http://www.msecm.com" name="MSECM(R) GmbH" phone="+49 8102 748397" state="BY" street="Ahornring 61" zip="85635"/></CONSTRUCTOR><MEETS><MEET city="Erlangen" course="LCM" deadline="2025-03-10" deadlinetime="19:00" hostclub="TB Erlangen" name="International Swim Meeting Erlangen 2025" nation="GER" organizer="TB Erlangen" timing="AUTOMATIC"><CONTACT city="Erlangen" country="GER" email="meldungen.schwimmen@tb-erlangen.de" name="Zebelein, Christian" phone="+49 176 32619612" street="Nägelsbachstr. 27" zip="91052"/><AGEDATE type="YEAR" value="2025-03-16"/><POOL name="Erlangen" lanemax="8" lanemin="1" type="INDOOR"/><POINTTABLE name="FINA Point Scoring Long Course 2023" version="2023"/><FEES/><QUALIFY conversion="NONE" from="2022-06-01" until="2023-05-01" percent="100"/><SESSIONS><SESSION course="LCM" date="2025-03-15" daytime="09:00" name="Abschnitt 1" number="1" warmupfrom="08:00" warmupuntil="09:00"><POOL name="Erlangen" lanemax="8" lanemin="1" type="INDOOR"/><JUDGES/><EVENTS><EVENT eventid="1" gender="F" number="1" order="1" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="700"/><SWIMSTYLE distance="50" name="50m Brust Frauen" relaycount="1" stroke="BREAST"/><AGEGROUPS><AGEGROUP agegroupid="10001" agemax="8" agemin="8" gender="F" name="Jahrgang 2017"><RANKINGS><RANKING place="5" resultid="7"/><RANKING place="6" resultid="8"/><RANKING place="2" resultid="16"/><RANKING place="8" resultid="20"/><RANKING place="3" resultid="25"/><RANKING place="7" resultid="28"/><RANKING place="4" resultid="36"/><RANKING place="-1" resultid="42"/><RANKING place="1" resultid="65"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="10002" agemax="9" agemin="9" gender="F" name="Jahrgang 2016"><RANKINGS><RANKING place="15" resultid="9"/><RANKING place="14" resultid="13"/><RANKING place="-1" resultid="19"/><RANKING place="13" resultid="21"/><RANKING place="5" resultid="22"/><RANKING place="11" resultid="24"/><RANKING place="12" resultid="26"/><RANKING place="4" resultid="31"/><RANKING place="7" resultid="33"/><RANKING place="10" resultid="38"/><RANKING place="6" resultid="43"/><RANKING place="9" resultid="45"/><RANKING place="8" resultid="51"/><RANKING place="2" resultid="57"/><RANKING place="3" resultid="60"/><RANKING place="1" resultid="95"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="10003" agemax="10" agemin="10" gender="F" name="Jahrgang 2015"><RANKINGS><RANKING place="26" resultid="2"/><RANKING place="24" resultid="11"/><RANKING place="25" resultid="12"/><RANKING place="21" resultid="29"/><RANKING place="18" resultid="30"/><RANKING place="13" resultid="32"/><RANKING place="20" resultid="37"/><RANKING place="19" resultid="40"/><RANKING place="14" resultid="41"/><RANKING place="16" resultid="47"/><RANKING place="17" resultid="48"/><RANKING place="15" resultid="49"/><RANKING place="-1" resultid="50"/><RANKING place="23" resultid="52"/><RANKING place="8" resultid="61"/><RANKING place="22" resultid="62"/><RANKING place="11" resultid="69"/><RANKING place="10" resultid="71"/><RANKING place="5" resultid="72"/><RANKING place="12" resultid="74"/><RANKING place="6" resultid="77"/><RANKING place="7" resultid="83"/><RANKING place="9" resultid="86"/><RANKING place="4" resultid="91"/><RANKING place="3" resultid="97"/><RANKING place="2" resultid="108"/><RANKING place="1" resultid="117"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="10004" agemax="11" agemin="11" gender="F" name="Jahrgang 2014"><RANKINGS><RANKING place="18" resultid="3"/><RANKING place="32" resultid="10"/><RANKING place="30" resultid="18"/><RANKING place="28" resultid="27"/><RANKING place="26" resultid="34"/><RANKING place="29" resultid="35"/><RANKING place="20" resultid="39"/><RANKING place="31" resultid="44"/><RANKING place="24" resultid="46"/><RANKING place="19" resultid="53"/><RANKING place="22" resultid="54"/><RANKING place="17" resultid="55"/><RANKING place="12" resultid="56"/><RANKING place="23" resultid="59"/><RANKING place="26" resultid="63"/><RANKING place="25" resultid="67"/><RANKING place="9" resultid="68"/><RANKING place="21" resultid="76"/><RANKING place="10" resultid="79"/><RANKING place="-1" resultid="80"/><RANKING place="15" resultid="82"/><RANKING place="14" resultid="84"/><RANKING place="-1" resultid="87"/><RANKING place="5" resultid="88"/><RANKING place="16" resultid="89"/><RANKING place="7" resultid="96"/><RANKING place="3" resultid="102"/><RANKING place="4" resultid="105"/><RANKING place="11" resultid="106"/><RANKING place="6" resultid="107"/><RANKING place="2" resultid="112"/><RANKING place="8" resultid="116"/><RANKING place="1" resultid="120"/><RANKING place="13" resultid="124"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="10005" agemax="12" agemin="12" gender="F" name="Jahrgang 2013"><RANKINGS><RANKING place="-1" resultid="1"/><RANKING place="19" resultid="6"/><RANKING place="-1" resultid="14"/><RANKING place="21" resultid="15"/><RANKING place="20" resultid="17"/><RANKING place="22" resultid="23"/><RANKING place="16" resultid="58"/><RANKING place="9" resultid="64"/><RANKING place="14" resultid="66"/><RANKING place="17" resultid="70"/><RANKING place="6" resultid="73"/><RANKING place="18" resultid="75"/><RANKING place="15" resultid="78"/><RANKING place="7" resultid="81"/><RANKING place="5" resultid="90"/><RANKING place="11" resultid="92"/><RANKING place="12" resultid="98"/><RANKING place="-1" resultid="101"/><RANKING place="8" resultid="103"/><RANKING place="10" resultid="110"/><RANKING place="2" resultid="114"/><RANKING place="13" resultid="115"/><RANKING place="-1" resultid="125"/><RANKING place="4" resultid="127"/><RANKING place="1" resultid="130"/><RANKING place="3" resultid="148"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="10006" agemax="13" agemin="13" gender="F" name="Jahrgang 2012"><RANKINGS><RANKING place="10" resultid="4"/><RANKING place="11" resultid="85"/><RANKING place="9" resultid="111"/><RANKING place="8" resultid="118"/><RANKING place="6" resultid="128"/><RANKING place="7" resultid="132"/><RANKING place="3" resultid="151"/><RANKING place="4" resultid="154"/><RANKING place="5" resultid="164"/><RANKING place="2" resultid="165"/><RANKING place="1" resultid="177"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="10007" agemax="14" agemin="14" gender="F" name="Jahrgang 2011"><RANKINGS><RANKING place="17" resultid="5"/><RANKING place="21" resultid="100"/><RANKING place="19" resultid="104"/><RANKING place="18" resultid="113"/><RANKING place="14" resultid="122"/><RANKING place="20" resultid="123"/><RANKING place="15" resultid="126"/><RANKING place="13" resultid="135"/><RANKING place="16" resultid="138"/><RANKING place="8" resultid="145"/><RANKING place="11" resultid="147"/><RANKING place="12" resultid="150"/><RANKING place="10" resultid="153"/><RANKING place="9" resultid="155"/><RANKING place="5" resultid="158"/><RANKING place="7" resultid="160"/><RANKING place="4" resultid="161"/><RANKING place="3" resultid="171"/><RANKING place="2" resultid="176"/><RANKING place="6" resultid="181"/><RANKING place="1" resultid="185"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="10008" agemax="15" agemin="15" gender="F" name="Jahrgang 2010"><RANKINGS><RANKING place="9" resultid="109"/><RANKING place="10" resultid="119"/><RANKING place="6" resultid="121"/><RANKING place="7" resultid="131"/><RANKING place="8" resultid="134"/><RANKING place="4" resultid="144"/><RANKING place="5" resultid="149"/><RANKING place="3" resultid="163"/><RANKING place="1" resultid="183"/><RANKING place="2" resultid="184"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="10009" agemax="16" agemin="16" gender="F" name="Jahrgang 2009"><RANKINGS><RANKING place="10" resultid="93"/><RANKING place="9" resultid="94"/><RANKING place="11" resultid="99"/><RANKING place="-1" resultid="129"/><RANKING place="-1" resultid="133"/><RANKING place="5" resultid="136"/><RANKING place="7" resultid="141"/><RANKING place="8" resultid="142"/><RANKING place="6" resultid="146"/><RANKING place="-1" resultid="166"/><RANKING place="4" resultid="168"/><RANKING place="2" resultid="169"/><RANKING place="3" resultid="172"/><RANKING place="1" resultid="173"/><RANKING place="-1" resultid="174"/><RANKING place="-1" resultid="179"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="10010" agemax="17" agemin="17" gender="F" name="Jahrgang 2008"><RANKINGS><RANKING place="2" resultid="143"/><RANKING place="1" resultid="159"/><RANKING place="-1" resultid="162"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="10011" agemax="-1" agemin="18" gender="F" name="Jahrgang 2007 und älter"><RANKINGS><RANKING place="13" resultid="137"/><RANKING place="11" resultid="139"/><RANKING place="9" resultid="140"/><RANKING place="6" resultid="152"/><RANKING place="8" resultid="156"/><RANKING place="12" resultid="157"/><RANKING place="4" resultid="167"/><RANKING place="10" resultid="170"/><RANKING place="2" resultid="175"/><RANKING place="7" resultid="178"/><RANKING place="3" resultid="180"/><RANKING place="1" resultid="182"/><RANKING place="5" resultid="186"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="1" number="1" order="1" status="OFFICIAL"/><HEAT heatid="2" number="2" order="2" status="OFFICIAL"/><HEAT heatid="3" number="3" order="3" status="OFFICIAL"/><HEAT heatid="4" number="4" order="4" status="OFFICIAL"/><HEAT heatid="5" number="5" order="5" status="OFFICIAL"/><HEAT heatid="6" number="6" order="6" status="OFFICIAL"/><HEAT heatid="7" number="7" order="7" status="OFFICIAL"/><HEAT heatid="8" number="8" order="8" status="OFFICIAL"/><HEAT heatid="9" number="9" order="9" status="OFFICIAL"/><HEAT heatid="10" number="10" order="10" status="OFFICIAL"/><HEAT heatid="11" number="11" order="11" status="OFFICIAL"/><HEAT heatid="12" number="12" order="12" status="OFFICIAL"/><HEAT heatid="13" number="13" order="13" status="OFFICIAL"/><HEAT heatid="14" number="14" order="14" status="OFFICIAL"/><HEAT heatid="15" number="15" order="15" status="OFFICIAL"/><HEAT heatid="16" number="16" order="16" status="OFFICIAL"/><HEAT heatid="17" number="17" order="17" status="OFFICIAL"/><HEAT heatid="18" number="18" order="18" status="OFFICIAL"/><HEAT heatid="19" number="19" order="19" status="OFFICIAL"/><HEAT heatid="20" number="20" order="20" status="OFFICIAL"/><HEAT heatid="21" number="21" order="21" status="OFFICIAL"/><HEAT heatid="22" number="22" order="22" status="OFFICIAL"/><HEAT heatid="23" number="23" order="23" status="OFFICIAL"/><HEAT heatid="24" number="24" order="24" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT><EVENT eventid="2" gender="M" number="2" order="2" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="700"/><SWIMSTYLE distance="50" name="50m Brust Männer" relaycount="1" stroke="BREAST"/><AGEGROUPS><AGEGROUP agegroupid="20001" agemax="8" agemin="8" gender="M" name="Jahrgang 2017"><RANKINGS><RANKING place="2" resultid="188"/><RANKING place="-1" resultid="189"/><RANKING place="1" resultid="204"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="20002" agemax="9" agemin="9" gender="M" name="Jahrgang 2016"><RANKINGS><RANKING place="7" resultid="190"/><RANKING place="-1" resultid="191"/><RANKING place="8" resultid="192"/><RANKING place="3" resultid="193"/><RANKING place="6" resultid="196"/><RANKING place="5" resultid="197"/><RANKING place="4" resultid="198"/><RANKING place="2" resultid="203"/><RANKING place="1" resultid="231"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="20003" agemax="10" agemin="10" gender="M" name="Jahrgang 2015"><RANKINGS><RANKING place="13" resultid="199"/><RANKING place="7" resultid="200"/><RANKING place="12" resultid="202"/><RANKING place="8" resultid="205"/><RANKING place="9" resultid="206"/><RANKING place="11" resultid="208"/><RANKING place="10" resultid="209"/><RANKING place="6" resultid="223"/><RANKING place="2" resultid="227"/><RANKING place="3" resultid="229"/><RANKING place="4" resultid="234"/><RANKING place="5" resultid="236"/><RANKING place="1" resultid="245"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="20004" agemax="11" agemin="11" gender="M" name="Jahrgang 2014"><RANKINGS><RANKING place="8" resultid="201"/><RANKING place="15" resultid="210"/><RANKING place="-1" resultid="212"/><RANKING place="17" resultid="213"/><RANKING place="6" resultid="214"/><RANKING place="13" resultid="215"/><RANKING place="4" resultid="216"/><RANKING place="12" resultid="219"/><RANKING place="16" resultid="220"/><RANKING place="14" resultid="222"/><RANKING place="11" resultid="224"/><RANKING place="10" resultid="225"/><RANKING place="5" resultid="226"/><RANKING place="7" resultid="230"/><RANKING place="1" resultid="232"/><RANKING place="2" resultid="233"/><RANKING place="3" resultid="242"/><RANKING place="9" resultid="244"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="20005" agemax="12" agemin="12" gender="M" name="Jahrgang 2013"><RANKINGS><RANKING place="12" resultid="187"/><RANKING place="11" resultid="194"/><RANKING place="13" resultid="211"/><RANKING place="-1" resultid="217"/><RANKING place="-1" resultid="218"/><RANKING place="9" resultid="221"/><RANKING place="10" resultid="235"/><RANKING place="6" resultid="246"/><RANKING place="4" resultid="249"/><RANKING place="3" resultid="250"/><RANKING place="5" resultid="251"/><RANKING place="8" resultid="252"/><RANKING place="7" resultid="253"/><RANKING place="-1" resultid="255"/><RANKING place="1" resultid="257"/><RANKING place="2" resultid="269"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="20006" agemax="13" agemin="13" gender="M" name="Jahrgang 2012"><RANKINGS><RANKING place="9" resultid="207"/><RANKING place="6" resultid="238"/><RANKING place="7" resultid="239"/><RANKING place="-1" resultid="240"/><RANKING place="2" resultid="243"/><RANKING place="8" resultid="247"/><RANKING place="4" resultid="259"/><RANKING place="5" resultid="260"/><RANKING place="3" resultid="261"/><RANKING place="1" resultid="272"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="20007" agemax="14" agemin="14" gender="M" name="Jahrgang 2011"><RANKINGS><RANKING place="14" resultid="254"/><RANKING place="13" resultid="256"/><RANKING place="10" resultid="258"/><RANKING place="8" resultid="263"/><RANKING place="5" resultid="264"/><RANKING place="12" resultid="265"/><RANKING place="11" resultid="266"/><RANKING place="7" resultid="270"/><RANKING place="4" resultid="271"/><RANKING place="6" resultid="273"/><RANKING place="9" resultid="274"/><RANKING place="-1" resultid="278"/><RANKING place="3" resultid="281"/><RANKING place="2" resultid="282"/><RANKING place="1" resultid="287"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="20008" agemax="15" agemin="15" gender="M" name="Jahrgang 2010"><RANKINGS><RANKING place="-1" resultid="228"/><RANKING place="10" resultid="241"/><RANKING place="9" resultid="248"/><RANKING place="11" resultid="267"/><RANKING place="8" resultid="268"/><RANKING place="4" resultid="275"/><RANKING place="3" resultid="285"/><RANKING place="2" resultid="286"/><RANKING place="5" resultid="288"/><RANKING place="7" resultid="290"/><RANKING place="6" resultid="291"/><RANKING place="1" resultid="297"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="20009" agemax="16" agemin="16" gender="M" name="Jahrgang 2009"><RANKINGS><RANKING place="4" resultid="262"/><RANKING place="5" resultid="276"/><RANKING place="6" resultid="277"/><RANKING place="2" resultid="295"/><RANKING place="1" resultid="302"/><RANKING place="3" resultid="304"/><RANKING place="-1" resultid="305"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="20010" agemax="17" agemin="17" gender="M" name="Jahrgang 2008"><RANKINGS><RANKING place="-1" resultid="237"/><RANKING place="3" resultid="283"/><RANKING place="2" resultid="289"/><RANKING place="1" resultid="299"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="20011" agemax="-1" agemin="18" gender="M" name="Jahrgang 2007 und älter"><RANKINGS><RANKING place="13" resultid="195"/><RANKING place="12" resultid="279"/><RANKING place="11" resultid="280"/><RANKING place="9" resultid="284"/><RANKING place="6" resultid="292"/><RANKING place="8" resultid="293"/><RANKING place="5" resultid="294"/><RANKING place="7" resultid="296"/><RANKING place="10" resultid="298"/><RANKING place="3" resultid="300"/><RANKING place="1" resultid="301"/><RANKING place="4" resultid="303"/><RANKING place="2" resultid="306"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="25" number="1" order="1" status="OFFICIAL"/><HEAT heatid="26" number="2" order="2" status="OFFICIAL"/><HEAT heatid="27" number="3" order="3" status="OFFICIAL"/><HEAT heatid="28" number="4" order="4" status="OFFICIAL"/><HEAT heatid="29" number="5" order="5" status="OFFICIAL"/><HEAT heatid="30" number="6" order="6" status="OFFICIAL"/><HEAT heatid="31" number="7" order="7" status="OFFICIAL"/><HEAT heatid="32" number="8" order="8" status="OFFICIAL"/><HEAT heatid="33" number="9" order="9" status="OFFICIAL"/><HEAT heatid="34" number="10" order="10" status="OFFICIAL"/><HEAT heatid="35" number="11" order="11" status="OFFICIAL"/><HEAT heatid="36" number="12" order="12" status="OFFICIAL"/><HEAT heatid="37" number="13" order="13" status="OFFICIAL"/><HEAT heatid="38" number="14" order="14" status="OFFICIAL"/><HEAT heatid="39" number="15" order="15" status="OFFICIAL"/><HEAT heatid="40" number="16" order="16" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT><EVENT eventid="3" gender="F" number="3" order="3" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="700"/><SWIMSTYLE distance="400" name="400m Freistil Frauen" relaycount="1" stroke="FREE"/><AGEGROUPS><AGEGROUP agegroupid="30001" agemax="10" agemin="10" gender="F" name="Jahrgang 2015"><RANKINGS><RANKING place="2" resultid="321"/><RANKING place="1" resultid="351"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="30002" agemax="11" agemin="11" gender="F" name="Jahrgang 2014"><RANKINGS><RANKING place="12" resultid="307"/><RANKING place="11" resultid="312"/><RANKING place="6" resultid="314"/><RANKING place="13" resultid="315"/><RANKING place="9" resultid="317"/><RANKING place="10" resultid="323"/><RANKING place="-1" resultid="327"/><RANKING place="8" resultid="330"/><RANKING place="2" resultid="331"/><RANKING place="5" resultid="335"/><RANKING place="4" resultid="336"/><RANKING place="7" resultid="338"/><RANKING place="1" resultid="349"/><RANKING place="3" resultid="350"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="30003" agemax="12" agemin="12" gender="F" name="Jahrgang 2013"><RANKINGS><RANKING place="12" resultid="308"/><RANKING place="13" resultid="309"/><RANKING place="14" resultid="310"/><RANKING place="-1" resultid="313"/><RANKING place="-1" resultid="316"/><RANKING place="11" resultid="318"/><RANKING place="-1" resultid="322"/><RANKING place="8" resultid="325"/><RANKING place="10" resultid="326"/><RANKING place="9" resultid="332"/><RANKING place="6" resultid="343"/><RANKING place="7" resultid="348"/><RANKING place="5" resultid="352"/><RANKING place="2" resultid="356"/><RANKING place="3" resultid="367"/><RANKING place="4" resultid="368"/><RANKING place="1" resultid="371"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="30004" agemax="13" agemin="13" gender="F" name="Jahrgang 2012"><RANKINGS><RANKING place="11" resultid="320"/><RANKING place="10" resultid="334"/><RANKING place="9" resultid="340"/><RANKING place="8" resultid="342"/><RANKING place="4" resultid="354"/><RANKING place="6" resultid="359"/><RANKING place="2" resultid="361"/><RANKING place="3" resultid="362"/><RANKING place="7" resultid="364"/><RANKING place="5" resultid="365"/><RANKING place="1" resultid="385"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="30005" agemax="14" agemin="14" gender="F" name="Jahrgang 2011"><RANKINGS><RANKING place="12" resultid="319"/><RANKING place="14" resultid="324"/><RANKING place="13" resultid="328"/><RANKING place="11" resultid="333"/><RANKING place="15" resultid="339"/><RANKING place="10" resultid="344"/><RANKING place="-1" resultid="345"/><RANKING place="9" resultid="346"/><RANKING place="8" resultid="357"/><RANKING place="7" resultid="360"/><RANKING place="6" resultid="369"/><RANKING place="5" resultid="372"/><RANKING place="4" resultid="377"/><RANKING place="3" resultid="379"/><RANKING place="2" resultid="386"/><RANKING place="1" resultid="397"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="30006" agemax="15" agemin="15" gender="F" name="Jahrgang 2010"><RANKINGS><RANKING place="14" resultid="311"/><RANKING place="12" resultid="329"/><RANKING place="9" resultid="337"/><RANKING place="13" resultid="341"/><RANKING place="11" resultid="358"/><RANKING place="8" resultid="363"/><RANKING place="10" resultid="366"/><RANKING place="7" resultid="370"/><RANKING place="5" resultid="378"/><RANKING place="6" resultid="381"/><RANKING place="4" resultid="383"/><RANKING place="3" resultid="391"/><RANKING place="1" resultid="393"/><RANKING place="2" resultid="395"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="30007" agemax="16" agemin="16" gender="F" name="Jahrgang 2009"><RANKINGS><RANKING place="5" resultid="353"/><RANKING place="7" resultid="355"/><RANKING place="9" resultid="373"/><RANKING place="8" resultid="374"/><RANKING place="10" resultid="375"/><RANKING place="4" resultid="376"/><RANKING place="6" resultid="380"/><RANKING place="3" resultid="382"/><RANKING place="1" resultid="384"/><RANKING place="2" resultid="390"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="30008" agemax="17" agemin="17" gender="F" name="Jahrgang 2008"><RANKINGS><RANKING place="2" resultid="387"/><RANKING place="1" resultid="394"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="30009" agemax="-1" agemin="18" gender="F" name="Jahrgang 2007 und älter"><RANKINGS><RANKING place="5" resultid="347"/><RANKING place="3" resultid="388"/><RANKING place="4" resultid="389"/><RANKING place="1" resultid="392"/><RANKING place="2" resultid="396"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="41" number="1" order="1" status="OFFICIAL"/><HEAT heatid="42" number="2" order="2" status="OFFICIAL"/><HEAT heatid="43" number="3" order="3" status="OFFICIAL"/><HEAT heatid="44" number="4" order="4" status="OFFICIAL"/><HEAT heatid="45" number="5" order="5" status="OFFICIAL"/><HEAT heatid="46" number="6" order="6" status="OFFICIAL"/><HEAT heatid="47" number="7" order="7" status="OFFICIAL"/><HEAT heatid="48" number="8" order="8" status="OFFICIAL"/><HEAT heatid="49" number="9" order="9" status="OFFICIAL"/><HEAT heatid="50" number="10" order="10" status="OFFICIAL"/><HEAT heatid="51" number="11" order="11" status="OFFICIAL"/><HEAT heatid="52" number="12" order="12" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT><EVENT eventid="4" gender="M" number="4" order="4" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="700"/><SWIMSTYLE distance="400" name="400m Freistil Männer" relaycount="1" stroke="FREE"/><AGEGROUPS><AGEGROUP agegroupid="40001" agemax="10" agemin="10" gender="M" name="Jahrgang 2015"><RANKINGS><RANKING place="10" resultid="404"/><RANKING place="5" resultid="405"/><RANKING place="9" resultid="406"/><RANKING place="3" resultid="407"/><RANKING place="6" resultid="408"/><RANKING place="8" resultid="409"/><RANKING place="2" resultid="412"/><RANKING place="7" resultid="417"/><RANKING place="4" resultid="419"/><RANKING place="1" resultid="426"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="40002" agemax="11" agemin="11" gender="M" name="Jahrgang 2014"><RANKINGS><RANKING place="6" resultid="398"/><RANKING place="7" resultid="400"/><RANKING place="8" resultid="402"/><RANKING place="5" resultid="403"/><RANKING place="4" resultid="415"/><RANKING place="3" resultid="416"/><RANKING place="1" resultid="427"/><RANKING place="2" resultid="433"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="40003" agemax="12" agemin="12" gender="M" name="Jahrgang 2013"><RANKINGS><RANKING place="12" resultid="399"/><RANKING place="10" resultid="410"/><RANKING place="8" resultid="413"/><RANKING place="11" resultid="414"/><RANKING place="4" resultid="418"/><RANKING place="5" resultid="421"/><RANKING place="7" resultid="422"/><RANKING place="6" resultid="423"/><RANKING place="9" resultid="425"/><RANKING place="3" resultid="436"/><RANKING place="-1" resultid="438"/><RANKING place="2" resultid="441"/><RANKING place="1" resultid="442"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="40004" agemax="13" agemin="13" gender="M" name="Jahrgang 2012"><RANKINGS><RANKING place="6" resultid="411"/><RANKING place="-1" resultid="431"/><RANKING place="5" resultid="432"/><RANKING place="2" resultid="439"/><RANKING place="3" resultid="440"/><RANKING place="1" resultid="443"/><RANKING place="4" resultid="446"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="40005" agemax="14" agemin="14" gender="M" name="Jahrgang 2011"><RANKINGS><RANKING place="-1" resultid="420"/><RANKING place="12" resultid="424"/><RANKING place="10" resultid="430"/><RANKING place="11" resultid="434"/><RANKING place="8" resultid="437"/><RANKING place="7" resultid="445"/><RANKING place="9" resultid="448"/><RANKING place="4" resultid="449"/><RANKING place="5" resultid="450"/><RANKING place="3" resultid="452"/><RANKING place="5" resultid="454"/><RANKING place="2" resultid="460"/><RANKING place="1" resultid="461"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="40006" agemax="15" agemin="15" gender="M" name="Jahrgang 2010"><RANKINGS><RANKING place="8" resultid="429"/><RANKING place="7" resultid="435"/><RANKING place="6" resultid="447"/><RANKING place="4" resultid="451"/><RANKING place="5" resultid="455"/><RANKING place="3" resultid="458"/><RANKING place="2" resultid="459"/><RANKING place="1" resultid="466"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="40007" agemax="16" agemin="16" gender="M" name="Jahrgang 2009"><RANKINGS><RANKING place="7" resultid="428"/><RANKING place="-1" resultid="444"/><RANKING place="5" resultid="453"/><RANKING place="6" resultid="456"/><RANKING place="2" resultid="462"/><RANKING place="4" resultid="465"/><RANKING place="3" resultid="467"/><RANKING place="1" resultid="468"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="40008" agemax="17" agemin="17" gender="M" name="Jahrgang 2008"><RANKINGS/></AGEGROUP><AGEGROUP agegroupid="40009" agemax="-1" agemin="18" gender="M" name="Jahrgang 2007 und älter"><RANKINGS><RANKING place="4" resultid="401"/><RANKING place="2" resultid="457"/><RANKING place="1" resultid="463"/><RANKING place="3" resultid="464"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="53" number="1" order="1" status="OFFICIAL"/><HEAT heatid="54" number="2" order="2" status="OFFICIAL"/><HEAT heatid="55" number="3" order="3" status="OFFICIAL"/><HEAT heatid="56" number="4" order="4" status="OFFICIAL"/><HEAT heatid="57" number="5" order="5" status="OFFICIAL"/><HEAT heatid="58" number="6" order="6" status="OFFICIAL"/><HEAT heatid="59" number="7" order="7" status="OFFICIAL"/><HEAT heatid="60" number="8" order="8" status="OFFICIAL"/><HEAT heatid="61" number="9" order="9" status="OFFICIAL"/><HEAT heatid="62" number="10" order="10" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT><EVENT eventid="5" gender="F" number="5" order="5" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="700"/><SWIMSTYLE distance="100" name="100m Schmetterling Frauen" relaycount="1" stroke="FLY"/><AGEGROUPS><AGEGROUP agegroupid="50001" agemax="10" agemin="10" gender="F" name="Jahrgang 2015"><RANKINGS><RANKING place="1" resultid="469"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="50002" agemax="11" agemin="11" gender="F" name="Jahrgang 2014"><RANKINGS><RANKING place="1" resultid="471"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="50003" agemax="12" agemin="12" gender="F" name="Jahrgang 2013"><RANKINGS><RANKING place="10" resultid="472"/><RANKING place="11" resultid="473"/><RANKING place="-1" resultid="475"/><RANKING place="9" resultid="476"/><RANKING place="8" resultid="477"/><RANKING place="6" resultid="484"/><RANKING place="3" resultid="486"/><RANKING place="7" resultid="487"/><RANKING place="2" resultid="489"/><RANKING place="4" resultid="497"/><RANKING place="5" resultid="502"/><RANKING place="1" resultid="511"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="50004" agemax="13" agemin="13" gender="F" name="Jahrgang 2012"><RANKINGS><RANKING place="10" resultid="474"/><RANKING place="7" resultid="478"/><RANKING place="9" resultid="480"/><RANKING place="8" resultid="482"/><RANKING place="6" resultid="490"/><RANKING place="4" resultid="504"/><RANKING place="3" resultid="510"/><RANKING place="5" resultid="512"/><RANKING place="1" resultid="523"/><RANKING place="2" resultid="527"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="50005" agemax="14" agemin="14" gender="F" name="Jahrgang 2011"><RANKINGS><RANKING place="9" resultid="470"/><RANKING place="8" resultid="479"/><RANKING place="7" resultid="485"/><RANKING place="10" resultid="488"/><RANKING place="6" resultid="494"/><RANKING place="2" resultid="507"/><RANKING place="5" resultid="509"/><RANKING place="3" resultid="517"/><RANKING place="-1" resultid="518"/><RANKING place="4" resultid="519"/><RANKING place="1" resultid="528"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="50006" agemax="15" agemin="15" gender="F" name="Jahrgang 2010"><RANKINGS><RANKING place="9" resultid="481"/><RANKING place="10" resultid="483"/><RANKING place="5" resultid="491"/><RANKING place="8" resultid="493"/><RANKING place="6" resultid="495"/><RANKING place="7" resultid="496"/><RANKING place="4" resultid="506"/><RANKING place="3" resultid="516"/><RANKING place="2" resultid="524"/><RANKING place="1" resultid="525"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="50007" agemax="16" agemin="16" gender="F" name="Jahrgang 2009"><RANKINGS><RANKING place="6" resultid="498"/><RANKING place="7" resultid="499"/><RANKING place="5" resultid="500"/><RANKING place="-1" resultid="513"/><RANKING place="4" resultid="514"/><RANKING place="3" resultid="515"/><RANKING place="2" resultid="529"/><RANKING place="1" resultid="533"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="50008" agemax="17" agemin="17" gender="F" name="Jahrgang 2008"><RANKINGS><RANKING place="6" resultid="501"/><RANKING place="5" resultid="505"/><RANKING place="4" resultid="520"/><RANKING place="3" resultid="526"/><RANKING place="1" resultid="534"/><RANKING place="2" resultid="535"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="50009" agemax="-1" agemin="18" gender="F" name="Jahrgang 2007 und älter"><RANKINGS><RANKING place="8" resultid="492"/><RANKING place="7" resultid="503"/><RANKING place="6" resultid="508"/><RANKING place="5" resultid="521"/><RANKING place="4" resultid="522"/><RANKING place="2" resultid="530"/><RANKING place="1" resultid="531"/><RANKING place="3" resultid="532"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="63" number="1" order="1" status="OFFICIAL"/><HEAT heatid="64" number="2" order="2" status="OFFICIAL"/><HEAT heatid="65" number="3" order="3" status="OFFICIAL"/><HEAT heatid="66" number="4" order="4" status="OFFICIAL"/><HEAT heatid="67" number="5" order="5" status="OFFICIAL"/><HEAT heatid="68" number="6" order="6" status="OFFICIAL"/><HEAT heatid="69" number="7" order="7" status="OFFICIAL"/><HEAT heatid="70" number="8" order="8" status="OFFICIAL"/><HEAT heatid="71" number="9" order="9" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT><EVENT eventid="6" gender="M" number="6" order="6" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="700"/><SWIMSTYLE distance="100" name="100m Schmetterling Männer" relaycount="1" stroke="FLY"/><AGEGROUPS><AGEGROUP agegroupid="60001" agemax="10" agemin="10" gender="M" name="Jahrgang 2015"><RANKINGS><RANKING place="1" resultid="544"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="60002" agemax="11" agemin="11" gender="M" name="Jahrgang 2014"><RANKINGS><RANKING place="2" resultid="536"/><RANKING place="1" resultid="537"/><RANKING place="3" resultid="538"/><RANKING place="4" resultid="543"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="60003" agemax="12" agemin="12" gender="M" name="Jahrgang 2013"><RANKINGS><RANKING place="5" resultid="539"/><RANKING place="4" resultid="540"/><RANKING place="3" resultid="542"/><RANKING place="1" resultid="558"/><RANKING place="2" resultid="559"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="60004" agemax="13" agemin="13" gender="M" name="Jahrgang 2012"><RANKINGS><RANKING place="3" resultid="545"/><RANKING place="2" resultid="547"/><RANKING place="6" resultid="554"/><RANKING place="5" resultid="556"/><RANKING place="4" resultid="566"/><RANKING place="1" resultid="567"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="60005" agemax="14" agemin="14" gender="M" name="Jahrgang 2011"><RANKINGS><RANKING place="6" resultid="546"/><RANKING place="5" resultid="548"/><RANKING place="9" resultid="549"/><RANKING place="7" resultid="550"/><RANKING place="8" resultid="555"/><RANKING place="-1" resultid="562"/><RANKING place="4" resultid="571"/><RANKING place="2" resultid="574"/><RANKING place="3" resultid="582"/><RANKING place="1" resultid="588"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="60006" agemax="15" agemin="15" gender="M" name="Jahrgang 2010"><RANKINGS><RANKING place="12" resultid="541"/><RANKING place="7" resultid="551"/><RANKING place="13" resultid="552"/><RANKING place="10" resultid="553"/><RANKING place="9" resultid="563"/><RANKING place="8" resultid="564"/><RANKING place="11" resultid="565"/><RANKING place="5" resultid="568"/><RANKING place="6" resultid="572"/><RANKING place="4" resultid="583"/><RANKING place="3" resultid="592"/><RANKING place="2" resultid="596"/><RANKING place="1" resultid="603"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="60007" agemax="16" agemin="16" gender="M" name="Jahrgang 2009"><RANKINGS><RANKING place="10" resultid="560"/><RANKING place="7" resultid="569"/><RANKING place="9" resultid="570"/><RANKING place="8" resultid="576"/><RANKING place="1" resultid="585"/><RANKING place="3" resultid="586"/><RANKING place="6" resultid="589"/><RANKING place="5" resultid="593"/><RANKING place="4" resultid="597"/><RANKING place="2" resultid="604"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="60008" agemax="17" agemin="17" gender="M" name="Jahrgang 2008"><RANKINGS><RANKING place="4" resultid="557"/><RANKING place="3" resultid="573"/><RANKING place="-1" resultid="595"/><RANKING place="2" resultid="600"/><RANKING place="1" resultid="601"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="60009" agemax="-1" agemin="18" gender="M" name="Jahrgang 2007 und älter"><RANKINGS><RANKING place="11" resultid="561"/><RANKING place="9" resultid="575"/><RANKING place="8" resultid="577"/><RANKING place="14" resultid="578"/><RANKING place="10" resultid="579"/><RANKING place="15" resultid="580"/><RANKING place="13" resultid="581"/><RANKING place="7" resultid="584"/><RANKING place="12" resultid="587"/><RANKING place="3" resultid="590"/><RANKING place="5" resultid="591"/><RANKING place="4" resultid="594"/><RANKING place="6" resultid="598"/><RANKING place="2" resultid="599"/><RANKING place="1" resultid="602"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="72" number="1" order="1" status="OFFICIAL"/><HEAT heatid="73" number="2" order="2" status="OFFICIAL"/><HEAT heatid="74" number="3" order="3" status="OFFICIAL"/><HEAT heatid="75" number="4" order="4" status="OFFICIAL"/><HEAT heatid="76" number="5" order="5" status="OFFICIAL"/><HEAT heatid="77" number="6" order="6" status="OFFICIAL"/><HEAT heatid="78" number="7" order="7" status="OFFICIAL"/><HEAT heatid="79" number="8" order="8" status="OFFICIAL"/><HEAT heatid="80" number="9" order="9" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT><EVENT eventid="7" gender="F" number="7" order="7" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="700"/><SWIMSTYLE distance="200" name="200m Brust Frauen" relaycount="1" stroke="BREAST"/><AGEGROUPS><AGEGROUP agegroupid="70001" agemax="10" agemin="10" gender="F" name="Jahrgang 2015"><RANKINGS><RANKING place="11" resultid="605"/><RANKING place="5" resultid="607"/><RANKING place="8" resultid="610"/><RANKING place="7" resultid="614"/><RANKING place="9" resultid="617"/><RANKING place="6" resultid="621"/><RANKING place="3" resultid="625"/><RANKING place="10" resultid="632"/><RANKING place="4" resultid="635"/><RANKING place="2" resultid="642"/><RANKING place="1" resultid="648"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="70002" agemax="11" agemin="11" gender="F" name="Jahrgang 2014"><RANKINGS><RANKING place="18" resultid="606"/><RANKING place="21" resultid="608"/><RANKING place="10" resultid="611"/><RANKING place="19" resultid="612"/><RANKING place="5" resultid="615"/><RANKING place="20" resultid="616"/><RANKING place="16" resultid="619"/><RANKING place="14" resultid="620"/><RANKING place="11" resultid="622"/><RANKING place="3" resultid="623"/><RANKING place="8" resultid="624"/><RANKING place="12" resultid="626"/><RANKING place="7" resultid="627"/><RANKING place="-1" resultid="628"/><RANKING place="17" resultid="630"/><RANKING place="9" resultid="633"/><RANKING place="13" resultid="634"/><RANKING place="-1" resultid="637"/><RANKING place="15" resultid="640"/><RANKING place="4" resultid="645"/><RANKING place="2" resultid="650"/><RANKING place="1" resultid="652"/><RANKING place="6" resultid="659"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="70003" agemax="12" agemin="12" gender="F" name="Jahrgang 2013"><RANKINGS><RANKING place="17" resultid="609"/><RANKING place="-1" resultid="613"/><RANKING place="18" resultid="618"/><RANKING place="10" resultid="629"/><RANKING place="15" resultid="636"/><RANKING place="14" resultid="638"/><RANKING place="12" resultid="639"/><RANKING place="16" resultid="641"/><RANKING place="11" resultid="643"/><RANKING place="-1" resultid="644"/><RANKING place="13" resultid="646"/><RANKING place="5" resultid="651"/><RANKING place="6" resultid="655"/><RANKING place="-1" resultid="656"/><RANKING place="9" resultid="657"/><RANKING place="7" resultid="658"/><RANKING place="8" resultid="660"/><RANKING place="4" resultid="661"/><RANKING place="2" resultid="668"/><RANKING place="3" resultid="669"/><RANKING place="1" resultid="679"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="70004" agemax="13" agemin="13" gender="F" name="Jahrgang 2012"><RANKINGS><RANKING place="6" resultid="631"/><RANKING place="3" resultid="649"/><RANKING place="5" resultid="665"/><RANKING place="4" resultid="672"/><RANKING place="2" resultid="678"/><RANKING place="1" resultid="681"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="70005" agemax="14" agemin="14" gender="F" name="Jahrgang 2011"><RANKINGS><RANKING place="8" resultid="647"/><RANKING place="6" resultid="654"/><RANKING place="7" resultid="663"/><RANKING place="-1" resultid="664"/><RANKING place="4" resultid="667"/><RANKING place="5" resultid="671"/><RANKING place="3" resultid="674"/><RANKING place="2" resultid="684"/><RANKING place="1" resultid="688"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="70006" agemax="15" agemin="15" gender="F" name="Jahrgang 2010"><RANKINGS><RANKING place="5" resultid="670"/><RANKING place="3" resultid="675"/><RANKING place="4" resultid="682"/><RANKING place="1" resultid="686"/><RANKING place="2" resultid="687"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="70007" agemax="16" agemin="16" gender="F" name="Jahrgang 2009"><RANKINGS><RANKING place="7" resultid="673"/><RANKING place="-1" resultid="676"/><RANKING place="4" resultid="677"/><RANKING place="-1" resultid="680"/><RANKING place="3" resultid="683"/><RANKING place="5" resultid="685"/><RANKING place="6" resultid="689"/><RANKING place="-1" resultid="690"/><RANKING place="1" resultid="692"/><RANKING place="2" resultid="696"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="70008" agemax="17" agemin="17" gender="F" name="Jahrgang 2008"><RANKINGS/></AGEGROUP><AGEGROUP agegroupid="70009" agemax="-1" agemin="18" gender="F" name="Jahrgang 2007 und älter"><RANKINGS><RANKING place="7" resultid="653"/><RANKING place="6" resultid="662"/><RANKING place="5" resultid="666"/><RANKING place="2" resultid="691"/><RANKING place="1" resultid="693"/><RANKING place="4" resultid="694"/><RANKING place="3" resultid="695"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="81" number="1" order="1" status="OFFICIAL"/><HEAT heatid="82" number="2" order="2" status="OFFICIAL"/><HEAT heatid="83" number="3" order="3" status="OFFICIAL"/><HEAT heatid="84" number="4" order="4" status="OFFICIAL"/><HEAT heatid="85" number="5" order="5" status="OFFICIAL"/><HEAT heatid="86" number="6" order="6" status="OFFICIAL"/><HEAT heatid="87" number="7" order="7" status="OFFICIAL"/><HEAT heatid="88" number="8" order="8" status="OFFICIAL"/><HEAT heatid="89" number="9" order="9" status="OFFICIAL"/><HEAT heatid="90" number="10" order="10" status="OFFICIAL"/><HEAT heatid="91" number="11" order="11" status="OFFICIAL"/><HEAT heatid="92" number="12" order="12" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT><EVENT eventid="8" gender="M" number="8" order="8" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="700"/><SWIMSTYLE distance="200" name="200m Brust Männer" relaycount="1" stroke="BREAST"/><AGEGROUPS><AGEGROUP agegroupid="80001" agemax="10" agemin="10" gender="M" name="Jahrgang 2015"><RANKINGS><RANKING place="4" resultid="700"/><RANKING place="7" resultid="702"/><RANKING place="6" resultid="708"/><RANKING place="2" resultid="712"/><RANKING place="3" resultid="716"/><RANKING place="5" resultid="723"/><RANKING place="1" resultid="725"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="80002" agemax="11" agemin="11" gender="M" name="Jahrgang 2014"><RANKINGS><RANKING place="11" resultid="698"/><RANKING place="5" resultid="699"/><RANKING place="7" resultid="701"/><RANKING place="6" resultid="703"/><RANKING place="12" resultid="705"/><RANKING place="-1" resultid="707"/><RANKING place="10" resultid="709"/><RANKING place="9" resultid="710"/><RANKING place="8" resultid="711"/><RANKING place="2" resultid="714"/><RANKING place="4" resultid="715"/><RANKING place="3" resultid="720"/><RANKING place="1" resultid="734"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="80003" agemax="12" agemin="12" gender="M" name="Jahrgang 2013"><RANKINGS><RANKING place="10" resultid="704"/><RANKING place="8" resultid="713"/><RANKING place="11" resultid="717"/><RANKING place="-1" resultid="719"/><RANKING place="4" resultid="722"/><RANKING place="9" resultid="726"/><RANKING place="3" resultid="728"/><RANKING place="7" resultid="731"/><RANKING place="6" resultid="733"/><RANKING place="5" resultid="735"/><RANKING place="2" resultid="738"/><RANKING place="1" resultid="746"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="80004" agemax="13" agemin="13" gender="M" name="Jahrgang 2012"><RANKINGS><RANKING place="5" resultid="718"/><RANKING place="4" resultid="724"/><RANKING place="3" resultid="729"/><RANKING place="1" resultid="742"/><RANKING place="2" resultid="745"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="80005" agemax="14" agemin="14" gender="M" name="Jahrgang 2011"><RANKINGS><RANKING place="7" resultid="721"/><RANKING place="4" resultid="727"/><RANKING place="8" resultid="730"/><RANKING place="9" resultid="732"/><RANKING place="5" resultid="736"/><RANKING place="6" resultid="739"/><RANKING place="10" resultid="740"/><RANKING place="2" resultid="749"/><RANKING place="1" resultid="750"/><RANKING place="-1" resultid="752"/><RANKING place="3" resultid="756"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="80006" agemax="15" agemin="15" gender="M" name="Jahrgang 2010"><RANKINGS><RANKING place="3" resultid="697"/><RANKING place="8" resultid="706"/><RANKING place="2" resultid="737"/><RANKING place="6" resultid="741"/><RANKING place="4" resultid="744"/><RANKING place="5" resultid="747"/><RANKING place="7" resultid="748"/><RANKING place="1" resultid="754"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="80007" agemax="16" agemin="16" gender="M" name="Jahrgang 2009"><RANKINGS><RANKING place="3" resultid="751"/><RANKING place="5" resultid="755"/><RANKING place="1" resultid="759"/><RANKING place="2" resultid="762"/><RANKING place="4" resultid="763"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="80008" agemax="17" agemin="17" gender="M" name="Jahrgang 2008"><RANKINGS><RANKING place="3" resultid="743"/><RANKING place="1" resultid="757"/><RANKING place="2" resultid="761"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="80009" agemax="-1" agemin="18" gender="M" name="Jahrgang 2007 und älter"><RANKINGS><RANKING place="3" resultid="753"/><RANKING place="2" resultid="758"/><RANKING place="1" resultid="760"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="93" number="1" order="1" status="OFFICIAL"/><HEAT heatid="94" number="2" order="2" status="OFFICIAL"/><HEAT heatid="95" number="3" order="3" status="OFFICIAL"/><HEAT heatid="96" number="4" order="4" status="OFFICIAL"/><HEAT heatid="97" number="5" order="5" status="OFFICIAL"/><HEAT heatid="98" number="6" order="6" status="OFFICIAL"/><HEAT heatid="99" number="7" order="7" status="OFFICIAL"/><HEAT heatid="100" number="8" order="8" status="OFFICIAL"/><HEAT heatid="101" number="9" order="9" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT></EVENTS></SESSION><SESSION course="LCM" date="2025-03-15" daytime="14:00" name="Abschnitt 2" number="2" warmupfrom="13:00" warmupuntil="14:00"><POOL name="Erlangen" lanemax="8" lanemin="1" type="INDOOR"/><JUDGES/><EVENTS><EVENT eventid="9" gender="F" number="9" order="9" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="700"/><SWIMSTYLE distance="50" name="50m Freistil Frauen" relaycount="1" stroke="FREE"/><AGEGROUPS><AGEGROUP agegroupid="90001" agemax="8" agemin="8" gender="F" name="Jahrgang 2017"><RANKINGS><RANKING place="8" resultid="770"/><RANKING place="7" resultid="777"/><RANKING place="6" resultid="779"/><RANKING place="4" resultid="782"/><RANKING place="2" resultid="783"/><RANKING place="5" resultid="786"/><RANKING place="1" resultid="794"/><RANKING place="3" resultid="809"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="90002" agemax="9" agemin="9" gender="F" name="Jahrgang 2016"><RANKINGS><RANKING place="13" resultid="772"/><RANKING place="12" resultid="773"/><RANKING place="16" resultid="774"/><RANKING place="14" resultid="775"/><RANKING place="10" resultid="780"/><RANKING place="15" resultid="784"/><RANKING place="11" resultid="788"/><RANKING place="-1" resultid="792"/><RANKING place="8" resultid="798"/><RANKING place="6" resultid="799"/><RANKING place="5" resultid="812"/><RANKING place="9" resultid="814"/><RANKING place="7" resultid="820"/><RANKING place="2" resultid="825"/><RANKING place="1" resultid="826"/><RANKING place="4" resultid="833"/><RANKING place="3" resultid="857"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="90003" agemax="10" agemin="10" gender="F" name="Jahrgang 2015"><RANKINGS><RANKING place="23" resultid="768"/><RANKING place="14" resultid="781"/><RANKING place="17" resultid="785"/><RANKING place="21" resultid="787"/><RANKING place="22" resultid="790"/><RANKING place="13" resultid="793"/><RANKING place="20" resultid="795"/><RANKING place="8" resultid="796"/><RANKING place="-1" resultid="800"/><RANKING place="18" resultid="801"/><RANKING place="19" resultid="802"/><RANKING place="10" resultid="803"/><RANKING place="12" resultid="815"/><RANKING place="15" resultid="817"/><RANKING place="5" resultid="821"/><RANKING place="11" resultid="822"/><RANKING place="16" resultid="824"/><RANKING place="6" resultid="829"/><RANKING place="7" resultid="830"/><RANKING place="3" resultid="835"/><RANKING place="9" resultid="837"/><RANKING place="4" resultid="844"/><RANKING place="2" resultid="853"/><RANKING place="1" resultid="860"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="90004" agemax="11" agemin="11" gender="F" name="Jahrgang 2014"><RANKINGS><RANKING place="20" resultid="764"/><RANKING place="27" resultid="767"/><RANKING place="18" resultid="804"/><RANKING place="19" resultid="805"/><RANKING place="21" resultid="806"/><RANKING place="23" resultid="807"/><RANKING place="25" resultid="808"/><RANKING place="26" resultid="810"/><RANKING place="22" resultid="811"/><RANKING place="24" resultid="816"/><RANKING place="-1" resultid="818"/><RANKING place="15" resultid="828"/><RANKING place="17" resultid="831"/><RANKING place="11" resultid="832"/><RANKING place="14" resultid="838"/><RANKING place="13" resultid="839"/><RANKING place="16" resultid="840"/><RANKING place="10" resultid="841"/><RANKING place="6" resultid="843"/><RANKING place="9" resultid="847"/><RANKING place="12" resultid="856"/><RANKING place="7" resultid="858"/><RANKING place="8" resultid="867"/><RANKING place="2" resultid="868"/><RANKING place="5" resultid="869"/><RANKING place="4" resultid="870"/><RANKING place="3" resultid="879"/><RANKING place="1" resultid="894"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="90005" agemax="12" agemin="12" gender="F" name="Jahrgang 2013"><RANKINGS><RANKING place="-1" resultid="766"/><RANKING place="-1" resultid="771"/><RANKING place="24" resultid="776"/><RANKING place="23" resultid="778"/><RANKING place="21" resultid="789"/><RANKING place="20" resultid="791"/><RANKING place="22" resultid="797"/><RANKING place="19" resultid="813"/><RANKING place="18" resultid="819"/><RANKING place="17" resultid="823"/><RANKING place="14" resultid="827"/><RANKING place="15" resultid="834"/><RANKING place="-1" resultid="836"/><RANKING place="16" resultid="848"/><RANKING place="6" resultid="851"/><RANKING place="-1" resultid="855"/><RANKING place="11" resultid="861"/><RANKING place="13" resultid="864"/><RANKING place="12" resultid="865"/><RANKING place="10" resultid="866"/><RANKING place="7" resultid="872"/><RANKING place="8" resultid="873"/><RANKING place="9" resultid="882"/><RANKING place="2" resultid="889"/><RANKING place="5" resultid="890"/><RANKING place="4" resultid="906"/><RANKING place="3" resultid="924"/><RANKING place="1" resultid="946"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="90006" agemax="13" agemin="13" gender="F" name="Jahrgang 2012"><RANKINGS><RANKING place="18" resultid="765"/><RANKING place="17" resultid="849"/><RANKING place="16" resultid="850"/><RANKING place="14" resultid="863"/><RANKING place="13" resultid="876"/><RANKING place="12" resultid="881"/><RANKING place="15" resultid="888"/><RANKING place="9" resultid="893"/><RANKING place="11" resultid="898"/><RANKING place="5" resultid="899"/><RANKING place="8" resultid="900"/><RANKING place="7" resultid="903"/><RANKING place="10" resultid="904"/><RANKING place="2" resultid="908"/><RANKING place="1" resultid="939"/><RANKING place="3" resultid="941"/><RANKING place="6" resultid="943"/><RANKING place="4" resultid="959"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="90007" agemax="14" agemin="14" gender="F" name="Jahrgang 2011"><RANKINGS><RANKING place="26" resultid="769"/><RANKING place="24" resultid="842"/><RANKING place="27" resultid="845"/><RANKING place="28" resultid="846"/><RANKING place="22" resultid="859"/><RANKING place="25" resultid="874"/><RANKING place="17" resultid="880"/><RANKING place="19" resultid="886"/><RANKING place="23" resultid="891"/><RANKING place="10" resultid="910"/><RANKING place="20" resultid="913"/><RANKING place="-1" resultid="914"/><RANKING place="18" resultid="915"/><RANKING place="14" resultid="922"/><RANKING place="13" resultid="925"/><RANKING place="4" resultid="930"/><RANKING place="21" resultid="935"/><RANKING place="-1" resultid="937"/><RANKING place="11" resultid="942"/><RANKING place="12" resultid="948"/><RANKING place="9" resultid="950"/><RANKING place="16" resultid="951"/><RANKING place="2" resultid="954"/><RANKING place="5" resultid="958"/><RANKING place="15" resultid="966"/><RANKING place="3" resultid="967"/><RANKING place="7" resultid="969"/><RANKING place="8" resultid="970"/><RANKING place="5" resultid="971"/><RANKING place="1" resultid="978"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="90008" agemax="15" agemin="15" gender="F" name="Jahrgang 2010"><RANKINGS><RANKING place="22" resultid="871"/><RANKING place="21" resultid="885"/><RANKING place="16" resultid="892"/><RANKING place="20" resultid="896"/><RANKING place="19" resultid="897"/><RANKING place="17" resultid="905"/><RANKING place="13" resultid="907"/><RANKING place="15" resultid="920"/><RANKING place="11" resultid="921"/><RANKING place="18" resultid="927"/><RANKING place="10" resultid="932"/><RANKING place="-1" resultid="933"/><RANKING place="13" resultid="934"/><RANKING place="9" resultid="936"/><RANKING place="12" resultid="944"/><RANKING place="6" resultid="947"/><RANKING place="8" resultid="955"/><RANKING place="5" resultid="962"/><RANKING place="7" resultid="975"/><RANKING place="4" resultid="981"/><RANKING place="3" resultid="986"/><RANKING place="2" resultid="987"/><RANKING place="1" resultid="991"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="90009" agemax="16" agemin="16" gender="F" name="Jahrgang 2009"><RANKINGS><RANKING place="23" resultid="854"/><RANKING place="22" resultid="862"/><RANKING place="-1" resultid="875"/><RANKING place="21" resultid="877"/><RANKING place="16" resultid="887"/><RANKING place="20" resultid="895"/><RANKING place="17" resultid="901"/><RANKING place="19" resultid="902"/><RANKING place="18" resultid="911"/><RANKING place="9" resultid="918"/><RANKING place="-1" resultid="923"/><RANKING place="12" resultid="931"/><RANKING place="-1" resultid="938"/><RANKING place="13" resultid="940"/><RANKING place="15" resultid="952"/><RANKING place="11" resultid="953"/><RANKING place="7" resultid="956"/><RANKING place="6" resultid="957"/><RANKING place="14" resultid="961"/><RANKING place="10" resultid="965"/><RANKING place="3" resultid="973"/><RANKING place="8" resultid="974"/><RANKING place="4" resultid="980"/><RANKING place="5" resultid="983"/><RANKING place="1" resultid="984"/><RANKING place="2" resultid="994"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="90010" agemax="17" agemin="17" gender="F" name="Jahrgang 2008"><RANKINGS><RANKING place="5" resultid="884"/><RANKING place="6" resultid="916"/><RANKING place="-1" resultid="919"/><RANKING place="4" resultid="964"/><RANKING place="3" resultid="968"/><RANKING place="2" resultid="977"/><RANKING place="1" resultid="995"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="90011" agemax="-1" agemin="18" gender="F" name="Jahrgang 2007 und älter"><RANKINGS><RANKING place="23" resultid="852"/><RANKING place="22" resultid="878"/><RANKING place="19" resultid="883"/><RANKING place="20" resultid="909"/><RANKING place="18" resultid="912"/><RANKING place="16" resultid="917"/><RANKING place="21" resultid="926"/><RANKING place="-1" resultid="928"/><RANKING place="17" resultid="929"/><RANKING place="14" resultid="945"/><RANKING place="12" resultid="949"/><RANKING place="13" resultid="960"/><RANKING place="9" resultid="963"/><RANKING place="7" resultid="972"/><RANKING place="8" resultid="976"/><RANKING place="10" resultid="979"/><RANKING place="11" resultid="982"/><RANKING place="4" resultid="985"/><RANKING place="1" resultid="988"/><RANKING place="15" resultid="989"/><RANKING place="5" resultid="990"/><RANKING place="2" resultid="992"/><RANKING place="3" resultid="993"/><RANKING place="6" resultid="996"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="102" number="1" order="1" status="OFFICIAL"/><HEAT heatid="103" number="2" order="2" status="OFFICIAL"/><HEAT heatid="104" number="3" order="3" status="OFFICIAL"/><HEAT heatid="105" number="4" order="4" status="OFFICIAL"/><HEAT heatid="106" number="5" order="5" status="OFFICIAL"/><HEAT heatid="107" number="6" order="6" status="OFFICIAL"/><HEAT heatid="108" number="7" order="7" status="OFFICIAL"/><HEAT heatid="109" number="8" order="8" status="OFFICIAL"/><HEAT heatid="110" number="9" order="9" status="OFFICIAL"/><HEAT heatid="111" number="10" order="10" status="OFFICIAL"/><HEAT heatid="112" number="11" order="11" status="OFFICIAL"/><HEAT heatid="113" number="12" order="12" status="OFFICIAL"/><HEAT heatid="114" number="13" order="13" status="OFFICIAL"/><HEAT heatid="115" number="14" order="14" status="OFFICIAL"/><HEAT heatid="116" number="15" order="15" status="OFFICIAL"/><HEAT heatid="117" number="16" order="16" status="OFFICIAL"/><HEAT heatid="118" number="17" order="17" status="OFFICIAL"/><HEAT heatid="119" number="18" order="18" status="OFFICIAL"/><HEAT heatid="120" number="19" order="19" status="OFFICIAL"/><HEAT heatid="121" number="20" order="20" status="OFFICIAL"/><HEAT heatid="122" number="21" order="21" status="OFFICIAL"/><HEAT heatid="123" number="22" order="22" status="OFFICIAL"/><HEAT heatid="124" number="23" order="23" status="OFFICIAL"/><HEAT heatid="125" number="24" order="24" status="OFFICIAL"/><HEAT heatid="126" number="25" order="25" status="OFFICIAL"/><HEAT heatid="127" number="26" order="26" status="OFFICIAL"/><HEAT heatid="128" number="27" order="27" status="OFFICIAL"/><HEAT heatid="129" number="28" order="28" status="OFFICIAL"/><HEAT heatid="130" number="29" order="29" status="OFFICIAL"/><HEAT heatid="131" number="30" order="30" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT><EVENT eventid="10" gender="M" number="10" order="10" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="700"/><SWIMSTYLE distance="50" name="50m Freistil Männer" relaycount="1" stroke="FREE"/><AGEGROUPS><AGEGROUP agegroupid="100001" agemax="8" agemin="8" gender="M" name="Jahrgang 2017"><RANKINGS><RANKING place="2" resultid="1004"/><RANKING place="1" resultid="1006"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="100002" agemax="9" agemin="9" gender="M" name="Jahrgang 2016"><RANKINGS><RANKING place="8" resultid="1001"/><RANKING place="5" resultid="1002"/><RANKING place="9" resultid="1003"/><RANKING place="3" resultid="1007"/><RANKING place="7" resultid="1012"/><RANKING place="4" resultid="1015"/><RANKING place="6" resultid="1020"/><RANKING place="2" resultid="1026"/><RANKING place="1" resultid="1048"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="100003" agemax="10" agemin="10" gender="M" name="Jahrgang 2015"><RANKINGS><RANKING place="14" resultid="1009"/><RANKING place="15" resultid="1010"/><RANKING place="11" resultid="1013"/><RANKING place="17" resultid="1014"/><RANKING place="12" resultid="1017"/><RANKING place="10" resultid="1018"/><RANKING place="16" resultid="1019"/><RANKING place="9" resultid="1021"/><RANKING place="7" resultid="1024"/><RANKING place="6" resultid="1027"/><RANKING place="13" resultid="1028"/><RANKING place="4" resultid="1039"/><RANKING place="5" resultid="1042"/><RANKING place="3" resultid="1054"/><RANKING place="1" resultid="1057"/><RANKING place="8" resultid="1059"/><RANKING place="2" resultid="1082"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="100004" agemax="11" agemin="11" gender="M" name="Jahrgang 2014"><RANKINGS><RANKING place="22" resultid="1011"/><RANKING place="15" resultid="1023"/><RANKING place="21" resultid="1025"/><RANKING place="16" resultid="1029"/><RANKING place="18" resultid="1030"/><RANKING place="13" resultid="1031"/><RANKING place="19" resultid="1032"/><RANKING place="12" resultid="1034"/><RANKING place="20" resultid="1035"/><RANKING place="17" resultid="1036"/><RANKING place="9" resultid="1043"/><RANKING place="8" resultid="1045"/><RANKING place="14" resultid="1046"/><RANKING place="10" resultid="1049"/><RANKING place="7" resultid="1052"/><RANKING place="-1" resultid="1053"/><RANKING place="6" resultid="1056"/><RANKING place="11" resultid="1058"/><RANKING place="1" resultid="1060"/><RANKING place="4" resultid="1066"/><RANKING place="5" resultid="1074"/><RANKING place="3" resultid="1081"/><RANKING place="2" resultid="1092"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="100005" agemax="12" agemin="12" gender="M" name="Jahrgang 2013"><RANKINGS><RANKING place="13" resultid="1000"/><RANKING place="16" resultid="1008"/><RANKING place="18" resultid="1022"/><RANKING place="14" resultid="1033"/><RANKING place="15" resultid="1037"/><RANKING place="-1" resultid="1038"/><RANKING place="9" resultid="1040"/><RANKING place="17" resultid="1044"/><RANKING place="6" resultid="1050"/><RANKING place="10" resultid="1055"/><RANKING place="3" resultid="1062"/><RANKING place="12" resultid="1063"/><RANKING place="-1" resultid="1064"/><RANKING place="11" resultid="1065"/><RANKING place="8" resultid="1069"/><RANKING place="4" resultid="1071"/><RANKING place="7" resultid="1073"/><RANKING place="5" resultid="1079"/><RANKING place="2" resultid="1086"/><RANKING place="1" resultid="1089"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="100006" agemax="13" agemin="13" gender="M" name="Jahrgang 2012"><RANKINGS><RANKING place="11" resultid="997"/><RANKING place="-1" resultid="998"/><RANKING place="12" resultid="1005"/><RANKING place="9" resultid="1047"/><RANKING place="10" resultid="1051"/><RANKING place="8" resultid="1061"/><RANKING place="-1" resultid="1075"/><RANKING place="4" resultid="1076"/><RANKING place="5" resultid="1080"/><RANKING place="2" resultid="1084"/><RANKING place="7" resultid="1085"/><RANKING place="6" resultid="1095"/><RANKING place="3" resultid="1112"/><RANKING place="1" resultid="1130"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="100007" agemax="14" agemin="14" gender="M" name="Jahrgang 2011"><RANKINGS><RANKING place="29" resultid="1041"/><RANKING place="28" resultid="1068"/><RANKING place="13" resultid="1070"/><RANKING place="-1" resultid="1072"/><RANKING place="23" resultid="1077"/><RANKING place="26" resultid="1083"/><RANKING place="25" resultid="1087"/><RANKING place="10" resultid="1088"/><RANKING place="20" resultid="1090"/><RANKING place="18" resultid="1093"/><RANKING place="21" resultid="1094"/><RANKING place="24" resultid="1096"/><RANKING place="27" resultid="1097"/><RANKING place="15" resultid="1098"/><RANKING place="14" resultid="1101"/><RANKING place="16" resultid="1102"/><RANKING place="17" resultid="1103"/><RANKING place="22" resultid="1106"/><RANKING place="11" resultid="1107"/><RANKING place="11" resultid="1110"/><RANKING place="19" resultid="1115"/><RANKING place="8" resultid="1118"/><RANKING place="9" resultid="1119"/><RANKING place="7" resultid="1128"/><RANKING place="4" resultid="1129"/><RANKING place="6" resultid="1132"/><RANKING place="5" resultid="1135"/><RANKING place="3" resultid="1153"/><RANKING place="1" resultid="1155"/><RANKING place="2" resultid="1160"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="100008" agemax="15" agemin="15" gender="M" name="Jahrgang 2010"><RANKINGS><RANKING place="22" resultid="999"/><RANKING place="23" resultid="1067"/><RANKING place="13" resultid="1091"/><RANKING place="17" resultid="1099"/><RANKING place="16" resultid="1100"/><RANKING place="18" resultid="1104"/><RANKING place="21" resultid="1105"/><RANKING place="8" resultid="1109"/><RANKING place="15" resultid="1111"/><RANKING place="20" resultid="1113"/><RANKING place="19" resultid="1114"/><RANKING place="14" resultid="1116"/><RANKING place="12" resultid="1120"/><RANKING place="10" resultid="1121"/><RANKING place="9" resultid="1123"/><RANKING place="11" resultid="1127"/><RANKING place="5" resultid="1131"/><RANKING place="5" resultid="1133"/><RANKING place="7" resultid="1134"/><RANKING place="4" resultid="1143"/><RANKING place="3" resultid="1165"/><RANKING place="2" resultid="1172"/><RANKING place="1" resultid="1188"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="100009" agemax="16" agemin="16" gender="M" name="Jahrgang 2009"><RANKINGS><RANKING place="19" resultid="1108"/><RANKING place="18" resultid="1117"/><RANKING place="17" resultid="1122"/><RANKING place="16" resultid="1125"/><RANKING place="9" resultid="1126"/><RANKING place="15" resultid="1137"/><RANKING place="14" resultid="1139"/><RANKING place="20" resultid="1140"/><RANKING place="10" resultid="1142"/><RANKING place="7" resultid="1154"/><RANKING place="11" resultid="1157"/><RANKING place="12" resultid="1158"/><RANKING place="13" resultid="1161"/><RANKING place="8" resultid="1164"/><RANKING place="6" resultid="1169"/><RANKING place="3" resultid="1171"/><RANKING place="2" resultid="1174"/><RANKING place="5" resultid="1182"/><RANKING place="1" resultid="1187"/><RANKING place="4" resultid="1191"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="100010" agemax="17" agemin="17" gender="M" name="Jahrgang 2008"><RANKINGS><RANKING place="7" resultid="1078"/><RANKING place="8" resultid="1124"/><RANKING place="6" resultid="1138"/><RANKING place="5" resultid="1151"/><RANKING place="-1" resultid="1156"/><RANKING place="-1" resultid="1168"/><RANKING place="-1" resultid="1170"/><RANKING place="3" resultid="1177"/><RANKING place="4" resultid="1184"/><RANKING place="2" resultid="1185"/><RANKING place="1" resultid="1190"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="100011" agemax="-1" agemin="18" gender="M" name="Jahrgang 2007 und älter"><RANKINGS><RANKING place="24" resultid="1016"/><RANKING place="22" resultid="1136"/><RANKING place="17" resultid="1141"/><RANKING place="21" resultid="1144"/><RANKING place="23" resultid="1145"/><RANKING place="20" resultid="1146"/><RANKING place="16" resultid="1147"/><RANKING place="-1" resultid="1148"/><RANKING place="10" resultid="1149"/><RANKING place="9" resultid="1150"/><RANKING place="19" resultid="1152"/><RANKING place="11" resultid="1159"/><RANKING place="14" resultid="1162"/><RANKING place="12" resultid="1163"/><RANKING place="13" resultid="1166"/><RANKING place="8" resultid="1167"/><RANKING place="7" resultid="1173"/><RANKING place="18" resultid="1175"/><RANKING place="6" resultid="1176"/><RANKING place="5" resultid="1178"/><RANKING place="-1" resultid="1179"/><RANKING place="4" resultid="1180"/><RANKING place="3" resultid="1181"/><RANKING place="15" resultid="1183"/><RANKING place="1" resultid="1186"/><RANKING place="2" resultid="1189"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="132" number="1" order="1" status="OFFICIAL"/><HEAT heatid="133" number="2" order="2" status="OFFICIAL"/><HEAT heatid="134" number="3" order="3" status="OFFICIAL"/><HEAT heatid="135" number="4" order="4" status="OFFICIAL"/><HEAT heatid="136" number="5" order="5" status="OFFICIAL"/><HEAT heatid="137" number="6" order="6" status="OFFICIAL"/><HEAT heatid="138" number="7" order="7" status="OFFICIAL"/><HEAT heatid="139" number="8" order="8" status="OFFICIAL"/><HEAT heatid="140" number="9" order="9" status="OFFICIAL"/><HEAT heatid="141" number="10" order="10" status="OFFICIAL"/><HEAT heatid="142" number="11" order="11" status="OFFICIAL"/><HEAT heatid="143" number="12" order="12" status="OFFICIAL"/><HEAT heatid="144" number="13" order="13" status="OFFICIAL"/><HEAT heatid="145" number="14" order="14" status="OFFICIAL"/><HEAT heatid="146" number="15" order="15" status="OFFICIAL"/><HEAT heatid="147" number="16" order="16" status="OFFICIAL"/><HEAT heatid="148" number="17" order="17" status="OFFICIAL"/><HEAT heatid="149" number="18" order="18" status="OFFICIAL"/><HEAT heatid="150" number="19" order="19" status="OFFICIAL"/><HEAT heatid="151" number="20" order="20" status="OFFICIAL"/><HEAT heatid="152" number="21" order="21" status="OFFICIAL"/><HEAT heatid="153" number="22" order="22" status="OFFICIAL"/><HEAT heatid="154" number="23" order="23" status="OFFICIAL"/><HEAT heatid="155" number="24" order="24" status="OFFICIAL"/><HEAT heatid="156" number="25" order="25" status="OFFICIAL"/><HEAT heatid="157" number="26" order="26" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT><EVENT eventid="11" gender="F" number="11" order="11" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="700"/><SWIMSTYLE distance="200" name="200m Lagen Frauen" relaycount="1" stroke="MEDLEY"/><AGEGROUPS><AGEGROUP agegroupid="110001" agemax="10" agemin="10" gender="F" name="Jahrgang 2015"><RANKINGS><RANKING place="5" resultid="1193"/><RANKING place="6" resultid="1194"/><RANKING place="4" resultid="1209"/><RANKING place="3" resultid="1215"/><RANKING place="2" resultid="1226"/><RANKING place="1" resultid="1232"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="110002" agemax="11" agemin="11" gender="F" name="Jahrgang 2014"><RANKINGS><RANKING place="14" resultid="1192"/><RANKING place="20" resultid="1195"/><RANKING place="12" resultid="1197"/><RANKING place="19" resultid="1199"/><RANKING place="17" resultid="1201"/><RANKING place="16" resultid="1203"/><RANKING place="18" resultid="1204"/><RANKING place="10" resultid="1205"/><RANKING place="15" resultid="1206"/><RANKING place="-1" resultid="1210"/><RANKING place="11" resultid="1216"/><RANKING place="13" resultid="1217"/><RANKING place="8" resultid="1220"/><RANKING place="4" resultid="1228"/><RANKING place="5" resultid="1233"/><RANKING place="9" resultid="1234"/><RANKING place="-1" resultid="1236"/><RANKING place="6" resultid="1237"/><RANKING place="-1" resultid="1238"/><RANKING place="7" resultid="1244"/><RANKING place="3" resultid="1245"/><RANKING place="2" resultid="1252"/><RANKING place="1" resultid="1282"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="110003" agemax="12" agemin="12" gender="F" name="Jahrgang 2013"><RANKINGS><RANKING place="27" resultid="1198"/><RANKING place="26" resultid="1200"/><RANKING place="28" resultid="1202"/><RANKING place="21" resultid="1208"/><RANKING place="25" resultid="1211"/><RANKING place="14" resultid="1212"/><RANKING place="20" resultid="1214"/><RANKING place="24" resultid="1218"/><RANKING place="22" resultid="1221"/><RANKING place="23" resultid="1222"/><RANKING place="18" resultid="1223"/><RANKING place="-1" resultid="1225"/><RANKING place="19" resultid="1230"/><RANKING place="16" resultid="1235"/><RANKING place="10" resultid="1240"/><RANKING place="15" resultid="1243"/><RANKING place="17" resultid="1250"/><RANKING place="13" resultid="1251"/><RANKING place="12" resultid="1255"/><RANKING place="8" resultid="1261"/><RANKING place="7" resultid="1263"/><RANKING place="9" resultid="1265"/><RANKING place="11" resultid="1266"/><RANKING place="6" resultid="1276"/><RANKING place="5" resultid="1277"/><RANKING place="3" resultid="1278"/><RANKING place="1" resultid="1289"/><RANKING place="4" resultid="1290"/><RANKING place="2" resultid="1295"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="110004" agemax="13" agemin="13" gender="F" name="Jahrgang 2012"><RANKINGS><RANKING place="14" resultid="1213"/><RANKING place="13" resultid="1227"/><RANKING place="12" resultid="1256"/><RANKING place="9" resultid="1262"/><RANKING place="8" resultid="1264"/><RANKING place="7" resultid="1268"/><RANKING place="10" resultid="1273"/><RANKING place="11" resultid="1274"/><RANKING place="5" resultid="1275"/><RANKING place="6" resultid="1279"/><RANKING place="3" resultid="1293"/><RANKING place="4" resultid="1299"/><RANKING place="2" resultid="1307"/><RANKING place="1" resultid="1311"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="110005" agemax="14" agemin="14" gender="F" name="Jahrgang 2011"><RANKINGS><RANKING place="15" resultid="1196"/><RANKING place="13" resultid="1207"/><RANKING place="12" resultid="1224"/><RANKING place="14" resultid="1229"/><RANKING place="11" resultid="1231"/><RANKING place="-1" resultid="1246"/><RANKING place="10" resultid="1247"/><RANKING place="9" resultid="1257"/><RANKING place="-1" resultid="1267"/><RANKING place="8" resultid="1272"/><RANKING place="5" resultid="1286"/><RANKING place="7" resultid="1287"/><RANKING place="6" resultid="1297"/><RANKING place="4" resultid="1301"/><RANKING place="3" resultid="1303"/><RANKING place="2" resultid="1314"/><RANKING place="1" resultid="1321"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="110006" agemax="15" agemin="15" gender="F" name="Jahrgang 2010"><RANKINGS><RANKING place="12" resultid="1219"/><RANKING place="8" resultid="1248"/><RANKING place="9" resultid="1249"/><RANKING place="10" resultid="1258"/><RANKING place="11" resultid="1260"/><RANKING place="7" resultid="1269"/><RANKING place="6" resultid="1285"/><RANKING place="4" resultid="1288"/><RANKING place="3" resultid="1292"/><RANKING place="-1" resultid="1296"/><RANKING place="5" resultid="1298"/><RANKING place="1" resultid="1320"/><RANKING place="2" resultid="1322"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="110007" agemax="16" agemin="16" gender="F" name="Jahrgang 2009"><RANKINGS><RANKING place="13" resultid="1239"/><RANKING place="12" resultid="1242"/><RANKING place="10" resultid="1253"/><RANKING place="11" resultid="1254"/><RANKING place="8" resultid="1271"/><RANKING place="9" resultid="1281"/><RANKING place="7" resultid="1283"/><RANKING place="6" resultid="1300"/><RANKING place="5" resultid="1304"/><RANKING place="-1" resultid="1305"/><RANKING place="4" resultid="1313"/><RANKING place="2" resultid="1316"/><RANKING place="3" resultid="1317"/><RANKING place="1" resultid="1318"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="110008" agemax="17" agemin="17" gender="F" name="Jahrgang 2008"><RANKINGS><RANKING place="4" resultid="1284"/><RANKING place="3" resultid="1302"/><RANKING place="2" resultid="1309"/><RANKING place="1" resultid="1310"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="110009" agemax="-1" agemin="18" gender="F" name="Jahrgang 2007 und älter"><RANKINGS><RANKING place="11" resultid="1241"/><RANKING place="9" resultid="1259"/><RANKING place="10" resultid="1270"/><RANKING place="8" resultid="1280"/><RANKING place="2" resultid="1291"/><RANKING place="3" resultid="1294"/><RANKING place="6" resultid="1306"/><RANKING place="5" resultid="1308"/><RANKING place="7" resultid="1312"/><RANKING place="4" resultid="1315"/><RANKING place="1" resultid="1319"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="158" number="1" order="1" status="OFFICIAL"/><HEAT heatid="159" number="2" order="2" status="OFFICIAL"/><HEAT heatid="160" number="3" order="3" status="OFFICIAL"/><HEAT heatid="161" number="4" order="4" status="OFFICIAL"/><HEAT heatid="162" number="5" order="5" status="OFFICIAL"/><HEAT heatid="163" number="6" order="6" status="OFFICIAL"/><HEAT heatid="164" number="7" order="7" status="OFFICIAL"/><HEAT heatid="165" number="8" order="8" status="OFFICIAL"/><HEAT heatid="166" number="9" order="9" status="OFFICIAL"/><HEAT heatid="167" number="10" order="10" status="OFFICIAL"/><HEAT heatid="168" number="11" order="11" status="OFFICIAL"/><HEAT heatid="169" number="12" order="12" status="OFFICIAL"/><HEAT heatid="170" number="13" order="13" status="OFFICIAL"/><HEAT heatid="171" number="14" order="14" status="OFFICIAL"/><HEAT heatid="172" number="15" order="15" status="OFFICIAL"/><HEAT heatid="173" number="16" order="16" status="OFFICIAL"/><HEAT heatid="174" number="17" order="17" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT><EVENT eventid="12" gender="M" number="12" order="12" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="700"/><SWIMSTYLE distance="200" name="200m Lagen Männer" relaycount="1" stroke="MEDLEY"/><AGEGROUPS><AGEGROUP agegroupid="120001" agemax="10" agemin="10" gender="M" name="Jahrgang 2015"><RANKINGS><RANKING place="7" resultid="1324"/><RANKING place="5" resultid="1325"/><RANKING place="8" resultid="1326"/><RANKING place="9" resultid="1329"/><RANKING place="4" resultid="1332"/><RANKING place="6" resultid="1333"/><RANKING place="3" resultid="1340"/><RANKING place="1" resultid="1346"/><RANKING place="2" resultid="1357"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="120002" agemax="11" agemin="11" gender="M" name="Jahrgang 2014"><RANKINGS><RANKING place="-1" resultid="1328"/><RANKING place="9" resultid="1330"/><RANKING place="10" resultid="1331"/><RANKING place="7" resultid="1335"/><RANKING place="8" resultid="1336"/><RANKING place="6" resultid="1338"/><RANKING place="11" resultid="1342"/><RANKING place="5" resultid="1347"/><RANKING place="-1" resultid="1348"/><RANKING place="3" resultid="1350"/><RANKING place="3" resultid="1352"/><RANKING place="2" resultid="1360"/><RANKING place="1" resultid="1383"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="120003" agemax="12" agemin="12" gender="M" name="Jahrgang 2013"><RANKINGS><RANKING place="16" resultid="1327"/><RANKING place="17" resultid="1334"/><RANKING place="14" resultid="1339"/><RANKING place="15" resultid="1341"/><RANKING place="13" resultid="1344"/><RANKING place="12" resultid="1345"/><RANKING place="11" resultid="1349"/><RANKING place="10" resultid="1354"/><RANKING place="9" resultid="1355"/><RANKING place="7" resultid="1356"/><RANKING place="8" resultid="1365"/><RANKING place="6" resultid="1367"/><RANKING place="5" resultid="1377"/><RANKING place="1" resultid="1382"/><RANKING place="3" resultid="1385"/><RANKING place="4" resultid="1387"/><RANKING place="2" resultid="1397"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="120004" agemax="13" agemin="13" gender="M" name="Jahrgang 2012"><RANKINGS><RANKING place="-1" resultid="1337"/><RANKING place="-1" resultid="1364"/><RANKING place="10" resultid="1371"/><RANKING place="9" resultid="1376"/><RANKING place="6" resultid="1380"/><RANKING place="7" resultid="1381"/><RANKING place="1" resultid="1386"/><RANKING place="8" resultid="1388"/><RANKING place="3" resultid="1389"/><RANKING place="4" resultid="1391"/><RANKING place="5" resultid="1394"/><RANKING place="2" resultid="1400"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="120005" agemax="14" agemin="14" gender="M" name="Jahrgang 2011"><RANKINGS><RANKING place="20" resultid="1343"/><RANKING place="17" resultid="1351"/><RANKING place="15" resultid="1353"/><RANKING place="19" resultid="1358"/><RANKING place="13" resultid="1359"/><RANKING place="14" resultid="1361"/><RANKING place="12" resultid="1363"/><RANKING place="8" resultid="1368"/><RANKING place="11" resultid="1369"/><RANKING place="16" resultid="1373"/><RANKING place="9" resultid="1375"/><RANKING place="10" resultid="1379"/><RANKING place="-1" resultid="1395"/><RANKING place="7" resultid="1401"/><RANKING place="3" resultid="1405"/><RANKING place="-1" resultid="1406"/><RANKING place="6" resultid="1411"/><RANKING place="5" resultid="1412"/><RANKING place="1" resultid="1413"/><RANKING place="18" resultid="1416"/><RANKING place="4" resultid="1418"/><RANKING place="2" resultid="1427"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="120006" agemax="15" agemin="15" gender="M" name="Jahrgang 2010"><RANKINGS><RANKING place="15" resultid="1362"/><RANKING place="18" resultid="1366"/><RANKING place="14" resultid="1370"/><RANKING place="17" resultid="1372"/><RANKING place="16" resultid="1374"/><RANKING place="13" resultid="1384"/><RANKING place="12" resultid="1390"/><RANKING place="7" resultid="1392"/><RANKING place="11" resultid="1393"/><RANKING place="9" resultid="1396"/><RANKING place="10" resultid="1402"/><RANKING place="8" resultid="1403"/><RANKING place="6" resultid="1404"/><RANKING place="4" resultid="1414"/><RANKING place="3" resultid="1421"/><RANKING place="5" resultid="1422"/><RANKING place="2" resultid="1428"/><RANKING place="1" resultid="1432"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="120007" agemax="16" agemin="16" gender="M" name="Jahrgang 2009"><RANKINGS><RANKING place="4" resultid="1378"/><RANKING place="2" resultid="1408"/><RANKING place="3" resultid="1409"/><RANKING place="1" resultid="1426"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="120008" agemax="17" agemin="17" gender="M" name="Jahrgang 2008"><RANKINGS><RANKING place="1" resultid="1399"/><RANKING place="-1" resultid="1407"/><RANKING place="-1" resultid="1420"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="120009" agemax="-1" agemin="18" gender="M" name="Jahrgang 2007 und älter"><RANKINGS><RANKING place="14" resultid="1323"/><RANKING place="13" resultid="1398"/><RANKING place="11" resultid="1410"/><RANKING place="8" resultid="1415"/><RANKING place="9" resultid="1417"/><RANKING place="10" resultid="1419"/><RANKING place="12" resultid="1423"/><RANKING place="6" resultid="1424"/><RANKING place="5" resultid="1425"/><RANKING place="4" resultid="1429"/><RANKING place="3" resultid="1430"/><RANKING place="1" resultid="1431"/><RANKING place="2" resultid="1433"/><RANKING place="7" resultid="1434"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="175" number="1" order="1" status="OFFICIAL"/><HEAT heatid="176" number="2" order="2" status="OFFICIAL"/><HEAT heatid="177" number="3" order="3" status="OFFICIAL"/><HEAT heatid="178" number="4" order="4" status="OFFICIAL"/><HEAT heatid="179" number="5" order="5" status="OFFICIAL"/><HEAT heatid="180" number="6" order="6" status="OFFICIAL"/><HEAT heatid="181" number="7" order="7" status="OFFICIAL"/><HEAT heatid="182" number="8" order="8" status="OFFICIAL"/><HEAT heatid="183" number="9" order="9" status="OFFICIAL"/><HEAT heatid="184" number="10" order="10" status="OFFICIAL"/><HEAT heatid="185" number="11" order="11" status="OFFICIAL"/><HEAT heatid="186" number="12" order="12" status="OFFICIAL"/><HEAT heatid="187" number="13" order="13" status="OFFICIAL"/><HEAT heatid="188" number="14" order="14" status="OFFICIAL"/><HEAT heatid="189" number="15" order="15" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT><EVENT eventid="13" gender="F" number="13" order="13" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="700"/><SWIMSTYLE distance="100" name="100m Rücken Frauen" relaycount="1" stroke="BACK"/><AGEGROUPS><AGEGROUP agegroupid="130001" agemax="8" agemin="8" gender="F" name="Jahrgang 2017"><RANKINGS><RANKING place="5" resultid="1436"/><RANKING place="2" resultid="1438"/><RANKING place="3" resultid="1449"/><RANKING place="1" resultid="1450"/><RANKING place="4" resultid="1453"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="130002" agemax="9" agemin="9" gender="F" name="Jahrgang 2016"><RANKINGS><RANKING place="10" resultid="1439"/><RANKING place="-1" resultid="1442"/><RANKING place="8" resultid="1448"/><RANKING place="9" resultid="1458"/><RANKING place="3" resultid="1459"/><RANKING place="6" resultid="1466"/><RANKING place="7" resultid="1468"/><RANKING place="1" resultid="1477"/><RANKING place="4" resultid="1480"/><RANKING place="2" resultid="1486"/><RANKING place="5" resultid="1487"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="130003" agemax="10" agemin="10" gender="F" name="Jahrgang 2015"><RANKINGS><RANKING place="17" resultid="1441"/><RANKING place="18" resultid="1446"/><RANKING place="14" resultid="1447"/><RANKING place="19" resultid="1451"/><RANKING place="-1" resultid="1452"/><RANKING place="20" resultid="1454"/><RANKING place="9" resultid="1460"/><RANKING place="12" resultid="1463"/><RANKING place="15" resultid="1467"/><RANKING place="8" resultid="1469"/><RANKING place="16" resultid="1470"/><RANKING place="13" resultid="1471"/><RANKING place="3" resultid="1473"/><RANKING place="11" resultid="1474"/><RANKING place="7" resultid="1478"/><RANKING place="10" resultid="1479"/><RANKING place="6" resultid="1485"/><RANKING place="4" resultid="1488"/><RANKING place="2" resultid="1492"/><RANKING place="5" resultid="1505"/><RANKING place="1" resultid="1519"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="130004" agemax="11" agemin="11" gender="F" name="Jahrgang 2014"><RANKINGS><RANKING place="25" resultid="1435"/><RANKING place="24" resultid="1437"/><RANKING place="22" resultid="1440"/><RANKING place="23" resultid="1443"/><RANKING place="21" resultid="1444"/><RANKING place="20" resultid="1455"/><RANKING place="16" resultid="1456"/><RANKING place="17" resultid="1457"/><RANKING place="-1" resultid="1462"/><RANKING place="18" resultid="1464"/><RANKING place="19" resultid="1465"/><RANKING place="14" resultid="1472"/><RANKING place="12" resultid="1475"/><RANKING place="-1" resultid="1476"/><RANKING place="11" resultid="1491"/><RANKING place="7" resultid="1493"/><RANKING place="15" resultid="1495"/><RANKING place="8" resultid="1496"/><RANKING place="9" resultid="1497"/><RANKING place="5" resultid="1499"/><RANKING place="6" resultid="1500"/><RANKING place="13" resultid="1503"/><RANKING place="4" resultid="1507"/><RANKING place="10" resultid="1510"/><RANKING place="2" resultid="1528"/><RANKING place="1" resultid="1538"/><RANKING place="3" resultid="1550"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="130005" agemax="12" agemin="12" gender="F" name="Jahrgang 2013"><RANKINGS><RANKING place="17" resultid="1445"/><RANKING place="16" resultid="1461"/><RANKING place="15" resultid="1484"/><RANKING place="13" resultid="1489"/><RANKING place="12" resultid="1490"/><RANKING place="9" resultid="1498"/><RANKING place="14" resultid="1501"/><RANKING place="10" resultid="1502"/><RANKING place="11" resultid="1506"/><RANKING place="-1" resultid="1509"/><RANKING place="7" resultid="1512"/><RANKING place="6" resultid="1520"/><RANKING place="8" resultid="1527"/><RANKING place="2" resultid="1530"/><RANKING place="4" resultid="1537"/><RANKING place="5" resultid="1544"/><RANKING place="1" resultid="1548"/><RANKING place="3" resultid="1573"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="130006" agemax="13" agemin="13" gender="F" name="Jahrgang 2012"><RANKINGS><RANKING place="8" resultid="1481"/><RANKING place="14" resultid="1482"/><RANKING place="13" resultid="1494"/><RANKING place="12" resultid="1511"/><RANKING place="11" resultid="1513"/><RANKING place="-1" resultid="1517"/><RANKING place="6" resultid="1523"/><RANKING place="7" resultid="1531"/><RANKING place="9" resultid="1532"/><RANKING place="4" resultid="1536"/><RANKING place="10" resultid="1541"/><RANKING place="5" resultid="1543"/><RANKING place="3" resultid="1545"/><RANKING place="2" resultid="1558"/><RANKING place="1" resultid="1588"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="130007" agemax="14" agemin="14" gender="F" name="Jahrgang 2011"><RANKINGS><RANKING place="16" resultid="1483"/><RANKING place="17" resultid="1508"/><RANKING place="13" resultid="1516"/><RANKING place="15" resultid="1521"/><RANKING place="-1" resultid="1525"/><RANKING place="12" resultid="1539"/><RANKING place="10" resultid="1546"/><RANKING place="5" resultid="1547"/><RANKING place="9" resultid="1551"/><RANKING place="8" resultid="1557"/><RANKING place="14" resultid="1560"/><RANKING place="3" resultid="1562"/><RANKING place="11" resultid="1564"/><RANKING place="7" resultid="1567"/><RANKING place="4" resultid="1570"/><RANKING place="6" resultid="1572"/><RANKING place="2" resultid="1582"/><RANKING place="1" resultid="1585"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="130008" agemax="15" agemin="15" gender="F" name="Jahrgang 2010"><RANKINGS><RANKING place="10" resultid="1504"/><RANKING place="7" resultid="1522"/><RANKING place="9" resultid="1535"/><RANKING place="8" resultid="1540"/><RANKING place="-1" resultid="1542"/><RANKING place="-1" resultid="1549"/><RANKING place="6" resultid="1552"/><RANKING place="4" resultid="1554"/><RANKING place="5" resultid="1559"/><RANKING place="3" resultid="1569"/><RANKING place="2" resultid="1576"/><RANKING place="1" resultid="1578"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="130009" agemax="16" agemin="16" gender="F" name="Jahrgang 2009"><RANKINGS><RANKING place="10" resultid="1514"/><RANKING place="12" resultid="1518"/><RANKING place="9" resultid="1529"/><RANKING place="11" resultid="1534"/><RANKING place="7" resultid="1555"/><RANKING place="8" resultid="1565"/><RANKING place="2" resultid="1579"/><RANKING place="5" resultid="1580"/><RANKING place="6" resultid="1581"/><RANKING place="3" resultid="1584"/><RANKING place="4" resultid="1586"/><RANKING place="1" resultid="1587"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="130010" agemax="17" agemin="17" gender="F" name="Jahrgang 2008"><RANKINGS><RANKING place="4" resultid="1515"/><RANKING place="5" resultid="1524"/><RANKING place="-1" resultid="1553"/><RANKING place="3" resultid="1561"/><RANKING place="2" resultid="1563"/><RANKING place="1" resultid="1571"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="130011" agemax="-1" agemin="18" gender="F" name="Jahrgang 2007 und älter"><RANKINGS><RANKING place="10" resultid="1526"/><RANKING place="9" resultid="1533"/><RANKING place="5" resultid="1556"/><RANKING place="7" resultid="1566"/><RANKING place="8" resultid="1568"/><RANKING place="6" resultid="1574"/><RANKING place="4" resultid="1575"/><RANKING place="3" resultid="1577"/><RANKING place="2" resultid="1583"/><RANKING place="1" resultid="1589"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="190" number="1" order="1" status="OFFICIAL"/><HEAT heatid="191" number="2" order="2" status="OFFICIAL"/><HEAT heatid="192" number="3" order="3" status="OFFICIAL"/><HEAT heatid="193" number="4" order="4" status="OFFICIAL"/><HEAT heatid="194" number="5" order="5" status="OFFICIAL"/><HEAT heatid="195" number="6" order="6" status="OFFICIAL"/><HEAT heatid="196" number="7" order="7" status="OFFICIAL"/><HEAT heatid="197" number="8" order="8" status="OFFICIAL"/><HEAT heatid="198" number="9" order="9" status="OFFICIAL"/><HEAT heatid="199" number="10" order="10" status="OFFICIAL"/><HEAT heatid="200" number="11" order="11" status="OFFICIAL"/><HEAT heatid="201" number="12" order="12" status="OFFICIAL"/><HEAT heatid="202" number="13" order="13" status="OFFICIAL"/><HEAT heatid="203" number="14" order="14" status="OFFICIAL"/><HEAT heatid="204" number="15" order="15" status="OFFICIAL"/><HEAT heatid="205" number="16" order="16" status="OFFICIAL"/><HEAT heatid="206" number="17" order="17" status="OFFICIAL"/><HEAT heatid="207" number="18" order="18" status="OFFICIAL"/><HEAT heatid="208" number="19" order="19" status="OFFICIAL"/><HEAT heatid="209" number="20" order="20" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT><EVENT eventid="14" gender="M" number="14" order="14" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="700"/><SWIMSTYLE distance="100" name="100m Rücken Männer" relaycount="1" stroke="BACK"/><AGEGROUPS><AGEGROUP agegroupid="140001" agemax="8" agemin="8" gender="M" name="Jahrgang 2017"><RANKINGS/></AGEGROUP><AGEGROUP agegroupid="140002" agemax="9" agemin="9" gender="M" name="Jahrgang 2016"><RANKINGS><RANKING place="2" resultid="1594"/><RANKING place="5" resultid="1595"/><RANKING place="6" resultid="1596"/><RANKING place="3" resultid="1602"/><RANKING place="4" resultid="1604"/><RANKING place="1" resultid="1650"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="140003" agemax="10" agemin="10" gender="M" name="Jahrgang 2015"><RANKINGS><RANKING place="19" resultid="1590"/><RANKING place="16" resultid="1592"/><RANKING place="14" resultid="1593"/><RANKING place="-1" resultid="1597"/><RANKING place="17" resultid="1601"/><RANKING place="10" resultid="1608"/><RANKING place="18" resultid="1612"/><RANKING place="11" resultid="1616"/><RANKING place="13" resultid="1618"/><RANKING place="4" resultid="1621"/><RANKING place="6" resultid="1623"/><RANKING place="8" resultid="1626"/><RANKING place="15" resultid="1627"/><RANKING place="12" resultid="1630"/><RANKING place="9" resultid="1642"/><RANKING place="2" resultid="1643"/><RANKING place="7" resultid="1644"/><RANKING place="5" resultid="1649"/><RANKING place="1" resultid="1655"/><RANKING place="3" resultid="1666"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="140004" agemax="11" agemin="11" gender="M" name="Jahrgang 2014"><RANKINGS><RANKING place="23" resultid="1598"/><RANKING place="-1" resultid="1599"/><RANKING place="21" resultid="1605"/><RANKING place="19" resultid="1606"/><RANKING place="20" resultid="1610"/><RANKING place="13" resultid="1614"/><RANKING place="22" resultid="1615"/><RANKING place="16" resultid="1617"/><RANKING place="17" resultid="1620"/><RANKING place="12" resultid="1625"/><RANKING place="15" resultid="1629"/><RANKING place="18" resultid="1631"/><RANKING place="11" resultid="1632"/><RANKING place="7" resultid="1633"/><RANKING place="9" resultid="1635"/><RANKING place="6" resultid="1637"/><RANKING place="8" resultid="1638"/><RANKING place="14" resultid="1639"/><RANKING place="10" resultid="1641"/><RANKING place="3" resultid="1646"/><RANKING place="4" resultid="1648"/><RANKING place="5" resultid="1651"/><RANKING place="2" resultid="1667"/><RANKING place="1" resultid="1671"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="140005" agemax="12" agemin="12" gender="M" name="Jahrgang 2013"><RANKINGS><RANKING place="15" resultid="1591"/><RANKING place="14" resultid="1600"/><RANKING place="13" resultid="1603"/><RANKING place="12" resultid="1607"/><RANKING place="3" resultid="1611"/><RANKING place="11" resultid="1613"/><RANKING place="10" resultid="1622"/><RANKING place="-1" resultid="1628"/><RANKING place="8" resultid="1634"/><RANKING place="5" resultid="1636"/><RANKING place="9" resultid="1640"/><RANKING place="7" resultid="1645"/><RANKING place="4" resultid="1656"/><RANKING place="-1" resultid="1658"/><RANKING place="6" resultid="1662"/><RANKING place="2" resultid="1669"/><RANKING place="1" resultid="1675"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="140006" agemax="13" agemin="13" gender="M" name="Jahrgang 2012"><RANKINGS><RANKING place="10" resultid="1609"/><RANKING place="9" resultid="1624"/><RANKING place="7" resultid="1653"/><RANKING place="5" resultid="1657"/><RANKING place="8" resultid="1659"/><RANKING place="6" resultid="1661"/><RANKING place="3" resultid="1670"/><RANKING place="4" resultid="1678"/><RANKING place="2" resultid="1688"/><RANKING place="1" resultid="1689"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="140007" agemax="14" agemin="14" gender="M" name="Jahrgang 2011"><RANKINGS><RANKING place="12" resultid="1619"/><RANKING place="11" resultid="1647"/><RANKING place="10" resultid="1652"/><RANKING place="7" resultid="1654"/><RANKING place="8" resultid="1660"/><RANKING place="5" resultid="1663"/><RANKING place="-1" resultid="1664"/><RANKING place="9" resultid="1665"/><RANKING place="6" resultid="1672"/><RANKING place="4" resultid="1673"/><RANKING place="-1" resultid="1679"/><RANKING place="3" resultid="1683"/><RANKING place="1" resultid="1684"/><RANKING place="2" resultid="1685"/><RANKING place="-1" resultid="1687"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="140008" agemax="15" agemin="15" gender="M" name="Jahrgang 2010"><RANKINGS><RANKING place="9" resultid="1668"/><RANKING place="7" resultid="1674"/><RANKING place="8" resultid="1680"/><RANKING place="6" resultid="1682"/><RANKING place="4" resultid="1686"/><RANKING place="5" resultid="1691"/><RANKING place="1" resultid="1699"/><RANKING place="2" resultid="1702"/><RANKING place="3" resultid="1704"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="140009" agemax="16" agemin="16" gender="M" name="Jahrgang 2009"><RANKINGS><RANKING place="8" resultid="1676"/><RANKING place="9" resultid="1681"/><RANKING place="6" resultid="1692"/><RANKING place="7" resultid="1696"/><RANKING place="4" resultid="1697"/><RANKING place="3" resultid="1698"/><RANKING place="5" resultid="1700"/><RANKING place="2" resultid="1701"/><RANKING place="1" resultid="1708"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="140010" agemax="17" agemin="17" gender="M" name="Jahrgang 2008"><RANKINGS><RANKING place="2" resultid="1690"/><RANKING place="-1" resultid="1695"/><RANKING place="-1" resultid="1703"/><RANKING place="1" resultid="1707"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="140011" agemax="-1" agemin="18" gender="M" name="Jahrgang 2007 und älter"><RANKINGS><RANKING place="6" resultid="1677"/><RANKING place="5" resultid="1693"/><RANKING place="-1" resultid="1694"/><RANKING place="3" resultid="1705"/><RANKING place="-1" resultid="1706"/><RANKING place="2" resultid="1709"/><RANKING place="1" resultid="1710"/><RANKING place="4" resultid="1711"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="210" number="1" order="1" status="OFFICIAL"/><HEAT heatid="211" number="2" order="2" status="OFFICIAL"/><HEAT heatid="212" number="3" order="3" status="OFFICIAL"/><HEAT heatid="213" number="4" order="4" status="OFFICIAL"/><HEAT heatid="214" number="5" order="5" status="OFFICIAL"/><HEAT heatid="215" number="6" order="6" status="OFFICIAL"/><HEAT heatid="216" number="7" order="7" status="OFFICIAL"/><HEAT heatid="217" number="8" order="8" status="OFFICIAL"/><HEAT heatid="218" number="9" order="9" status="OFFICIAL"/><HEAT heatid="219" number="10" order="10" status="OFFICIAL"/><HEAT heatid="220" number="11" order="11" status="OFFICIAL"/><HEAT heatid="221" number="12" order="12" status="OFFICIAL"/><HEAT heatid="222" number="13" order="13" status="OFFICIAL"/><HEAT heatid="223" number="14" order="14" status="OFFICIAL"/><HEAT heatid="224" number="15" order="15" status="OFFICIAL"/><HEAT heatid="225" number="16" order="16" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT></EVENTS></SESSION><SESSION course="LCM" date="2025-03-15" daytime="18:15" name="Abschnitt 3" number="3" warmupfrom="18:00" warmupuntil="18:15"><POOL name="Erlangen" lanemax="8" lanemin="1" type="INDOOR"/><JUDGES/><EVENTS><EVENT eventid="15" gender="F" number="15" order="15" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="1500"/><SWIMSTYLE distance="1500" name="1500m Freistil Frauen" relaycount="1" stroke="FREE"/><AGEGROUPS><AGEGROUP agegroupid="150001" agemax="-1" agemin="11" gender="F" name="Jahrgang 2014 und älter"><RANKINGS><RANKING place="10" resultid="1712"/><RANKING place="9" resultid="1713"/><RANKING place="8" resultid="1714"/><RANKING place="11" resultid="1715"/><RANKING place="5" resultid="1716"/><RANKING place="7" resultid="1717"/><RANKING place="4" resultid="1718"/><RANKING place="1" resultid="1719"/><RANKING place="2" resultid="1720"/><RANKING place="6" resultid="1721"/><RANKING place="3" resultid="1722"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="226" number="1" order="1" status="OFFICIAL"/><HEAT heatid="227" number="2" order="2" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT><EVENT eventid="16" gender="M" number="16" order="16" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="1500"/><SWIMSTYLE distance="1500" name="1500m Freistil Männer" relaycount="1" stroke="FREE"/><AGEGROUPS><AGEGROUP agegroupid="160001" agemax="-1" agemin="11" gender="M" name="Jahrgang 2014 und älter"><RANKINGS><RANKING place="9" resultid="1723"/><RANKING place="6" resultid="1724"/><RANKING place="7" resultid="1725"/><RANKING place="5" resultid="1726"/><RANKING place="1" resultid="1727"/><RANKING place="8" resultid="1728"/><RANKING place="2" resultid="1729"/><RANKING place="3" resultid="1730"/><RANKING place="4" resultid="1731"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="228" number="1" order="1" status="OFFICIAL"/><HEAT heatid="229" number="2" order="2" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT><EVENT eventid="17" gender="F" number="17" order="17" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="1500"/><SWIMSTYLE distance="800" name="800m Freistil Frauen" relaycount="1" stroke="FREE"/><AGEGROUPS><AGEGROUP agegroupid="170001" agemax="-1" agemin="11" gender="F" name="Jahrgang 2014 und älter"><RANKINGS><RANKING place="11" resultid="1732"/><RANKING place="14" resultid="1733"/><RANKING place="8" resultid="1734"/><RANKING place="10" resultid="1735"/><RANKING place="9" resultid="1736"/><RANKING place="12" resultid="1737"/><RANKING place="-1" resultid="1738"/><RANKING place="15" resultid="1739"/><RANKING place="5" resultid="1740"/><RANKING place="4" resultid="1741"/><RANKING place="3" resultid="1742"/><RANKING place="1" resultid="1743"/><RANKING place="2" resultid="1744"/><RANKING place="13" resultid="1745"/><RANKING place="7" resultid="1746"/><RANKING place="6" resultid="1747"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="230" number="1" order="1" status="OFFICIAL"/><HEAT heatid="231" number="2" order="2" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT><EVENT eventid="18" gender="M" number="18" order="18" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="1500"/><SWIMSTYLE distance="800" name="800m Freistil Männer" relaycount="1" stroke="FREE"/><AGEGROUPS><AGEGROUP agegroupid="180001" agemax="-1" agemin="11" gender="M" name="Jahrgang 2014 und älter"><RANKINGS><RANKING place="10" resultid="1748"/><RANKING place="-1" resultid="1749"/><RANKING place="6" resultid="1750"/><RANKING place="3" resultid="1751"/><RANKING place="9" resultid="1752"/><RANKING place="8" resultid="1753"/><RANKING place="5" resultid="1754"/><RANKING place="2" resultid="1755"/><RANKING place="4" resultid="1756"/><RANKING place="1" resultid="1757"/><RANKING place="7" resultid="1758"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="232" number="1" order="1" status="OFFICIAL"/><HEAT heatid="233" number="2" order="2" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT></EVENTS></SESSION><SESSION course="LCM" date="2025-03-16" daytime="08:30" name="Abschnitt 4" number="4" warmupfrom="07:30" warmupuntil="08:30"><POOL name="Erlangen" lanemax="8" lanemin="1" type="INDOOR"/><JUDGES/><EVENTS><EVENT eventid="19" gender="F" number="19" order="19" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="700"/><SWIMSTYLE distance="50" name="50m Rücken Beine Frauen" relaycount="1" stroke="UNKNOWN" technique="KICK"/><AGEGROUPS><AGEGROUP agegroupid="190001" agemax="11" agemin="11" gender="F" name="Jahrgang 2014"><RANKINGS><RANKING place="6" resultid="1759"/><RANKING place="5" resultid="1762"/><RANKING place="2" resultid="1763"/><RANKING place="4" resultid="1764"/><RANKING place="3" resultid="1765"/><RANKING place="1" resultid="1768"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="190002" agemax="12" agemin="12" gender="F" name="Jahrgang 2013"><RANKINGS><RANKING place="3" resultid="1760"/><RANKING place="1" resultid="1761"/><RANKING place="-1" resultid="1766"/><RANKING place="2" resultid="1767"/><RANKING place="4" resultid="1769"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="234" number="1" order="1" status="OFFICIAL"/><HEAT heatid="235" number="2" order="2" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT><EVENT eventid="20" gender="M" number="20" order="20" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="700"/><SWIMSTYLE distance="50" name="50m Rücken Beine Männer" relaycount="1" stroke="UNKNOWN" technique="KICK"/><AGEGROUPS><AGEGROUP agegroupid="200001" agemax="11" agemin="11" gender="M" name="Jahrgang 2014"><RANKINGS><RANKING place="3" resultid="1770"/><RANKING place="2" resultid="1772"/><RANKING place="1" resultid="1773"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="200002" agemax="12" agemin="12" gender="M" name="Jahrgang 2013"><RANKINGS><RANKING place="2" resultid="1771"/><RANKING place="1" resultid="1774"/><RANKING place="3" resultid="1775"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="236" number="1" order="1" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT><EVENT eventid="21" gender="F" number="21" order="21" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="700"/><SWIMSTYLE distance="50" name="50m Schmetterling Beine Frauen" relaycount="1" stroke="UNKNOWN" technique="KICK"/><AGEGROUPS><AGEGROUP agegroupid="210001" agemax="11" agemin="11" gender="F" name="Jahrgang 2014"><RANKINGS><RANKING place="2" resultid="1776"/><RANKING place="1" resultid="1780"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="210002" agemax="12" agemin="12" gender="F" name="Jahrgang 2013"><RANKINGS><RANKING place="3" resultid="1777"/><RANKING place="4" resultid="1778"/><RANKING place="5" resultid="1779"/><RANKING place="-1" resultid="1781"/><RANKING place="2" resultid="1782"/><RANKING place="1" resultid="1783"/><RANKING place="6" resultid="1784"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="237" number="1" order="1" status="OFFICIAL"/><HEAT heatid="238" number="2" order="2" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT><EVENT eventid="22" gender="M" number="22" order="22" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="700"/><SWIMSTYLE distance="50" name="50m Schmetterling Beine Männer" relaycount="1" stroke="UNKNOWN" technique="KICK"/><AGEGROUPS><AGEGROUP agegroupid="220001" agemax="11" agemin="11" gender="M" name="Jahrgang 2014"><RANKINGS><RANKING place="3" resultid="1785"/><RANKING place="2" resultid="1788"/><RANKING place="1" resultid="1789"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="220002" agemax="12" agemin="12" gender="M" name="Jahrgang 2013"><RANKINGS><RANKING place="2" resultid="1786"/><RANKING place="1" resultid="1787"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="239" number="1" order="1" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT><EVENT eventid="23" gender="F" number="23" order="23" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="700"/><SWIMSTYLE distance="50" name="50m Freistil Beine Frauen" relaycount="1" stroke="UNKNOWN" technique="KICK"/><AGEGROUPS><AGEGROUP agegroupid="230001" agemax="11" agemin="11" gender="F" name="Jahrgang 2014"><RANKINGS><RANKING place="13" resultid="1790"/><RANKING place="9" resultid="1792"/><RANKING place="6" resultid="1794"/><RANKING place="8" resultid="1797"/><RANKING place="12" resultid="1798"/><RANKING place="-1" resultid="1801"/><RANKING place="5" resultid="1802"/><RANKING place="10" resultid="1803"/><RANKING place="11" resultid="1804"/><RANKING place="2" resultid="1808"/><RANKING place="1" resultid="1809"/><RANKING place="7" resultid="1812"/><RANKING place="4" resultid="1813"/><RANKING place="3" resultid="1814"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="230002" agemax="12" agemin="12" gender="F" name="Jahrgang 2013"><RANKINGS><RANKING place="10" resultid="1791"/><RANKING place="2" resultid="1793"/><RANKING place="7" resultid="1795"/><RANKING place="8" resultid="1796"/><RANKING place="6" resultid="1799"/><RANKING place="5" resultid="1800"/><RANKING place="3" resultid="1805"/><RANKING place="9" resultid="1806"/><RANKING place="-1" resultid="1807"/><RANKING place="1" resultid="1810"/><RANKING place="4" resultid="1811"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="240" number="1" order="1" status="OFFICIAL"/><HEAT heatid="241" number="2" order="2" status="OFFICIAL"/><HEAT heatid="242" number="3" order="3" status="OFFICIAL"/><HEAT heatid="243" number="4" order="4" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT><EVENT eventid="24" gender="M" number="24" order="24" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="700"/><SWIMSTYLE distance="50" name="50m Freistil Beine Männer" relaycount="1" stroke="UNKNOWN" technique="KICK"/><AGEGROUPS><AGEGROUP agegroupid="240001" agemax="11" agemin="11" gender="M" name="Jahrgang 2014"><RANKINGS><RANKING place="3" resultid="1815"/><RANKING place="4" resultid="1818"/><RANKING place="2" resultid="1819"/><RANKING place="-1" resultid="1822"/><RANKING place="1" resultid="1824"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="240002" agemax="12" agemin="12" gender="M" name="Jahrgang 2013"><RANKINGS><RANKING place="8" resultid="1816"/><RANKING place="3" resultid="1817"/><RANKING place="6" resultid="1820"/><RANKING place="7" resultid="1821"/><RANKING place="2" resultid="1823"/><RANKING place="1" resultid="1825"/><RANKING place="5" resultid="1826"/><RANKING place="4" resultid="1827"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="244" number="1" order="1" status="OFFICIAL"/><HEAT heatid="245" number="2" order="2" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT><EVENT eventid="25" gender="F" number="25" order="25" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="700"/><SWIMSTYLE distance="50" name="50m Brust Beine Frauen" relaycount="1" stroke="UNKNOWN" technique="KICK"/><AGEGROUPS><AGEGROUP agegroupid="250001" agemax="11" agemin="11" gender="F" name="Jahrgang 2014"><RANKINGS><RANKING place="12" resultid="1828"/><RANKING place="8" resultid="1830"/><RANKING place="6" resultid="1833"/><RANKING place="7" resultid="1834"/><RANKING place="4" resultid="1837"/><RANKING place="3" resultid="1839"/><RANKING place="9" resultid="1842"/><RANKING place="11" resultid="1844"/><RANKING place="-1" resultid="1847"/><RANKING place="1" resultid="1848"/><RANKING place="5" resultid="1849"/><RANKING place="2" resultid="1850"/><RANKING place="10" resultid="1851"/><RANKING place="-1" resultid="1852"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="250002" agemax="12" agemin="12" gender="F" name="Jahrgang 2013"><RANKINGS><RANKING place="9" resultid="1829"/><RANKING place="3" resultid="1831"/><RANKING place="7" resultid="1832"/><RANKING place="6" resultid="1835"/><RANKING place="8" resultid="1836"/><RANKING place="-1" resultid="1838"/><RANKING place="1" resultid="1840"/><RANKING place="4" resultid="1841"/><RANKING place="2" resultid="1843"/><RANKING place="5" resultid="1845"/><RANKING place="-1" resultid="1846"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="246" number="1" order="1" status="OFFICIAL"/><HEAT heatid="247" number="2" order="2" status="OFFICIAL"/><HEAT heatid="248" number="3" order="3" status="OFFICIAL"/><HEAT heatid="249" number="4" order="4" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT><EVENT eventid="26" gender="M" number="26" order="26" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="700"/><SWIMSTYLE distance="50" name="50m Brust Beine Männer" relaycount="1" stroke="UNKNOWN" technique="KICK"/><AGEGROUPS><AGEGROUP agegroupid="260001" agemax="11" agemin="11" gender="M" name="Jahrgang 2014"><RANKINGS><RANKING place="5" resultid="1853"/><RANKING place="3" resultid="1854"/><RANKING place="1" resultid="1857"/><RANKING place="2" resultid="1860"/><RANKING place="4" resultid="1861"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="260002" agemax="12" agemin="12" gender="M" name="Jahrgang 2013"><RANKINGS><RANKING place="3" resultid="1855"/><RANKING place="2" resultid="1856"/><RANKING place="-1" resultid="1858"/><RANKING place="1" resultid="1859"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="250" number="1" order="1" status="OFFICIAL"/><HEAT heatid="251" number="2" order="2" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT><EVENT eventid="27" gender="F" number="27" order="27" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="700"/><SWIMSTYLE distance="50" name="50m Rücken Frauen" relaycount="1" stroke="BACK"/><AGEGROUPS><AGEGROUP agegroupid="270001" agemax="8" agemin="8" gender="F" name="Jahrgang 2017"><RANKINGS><RANKING place="7" resultid="1868"/><RANKING place="8" resultid="1874"/><RANKING place="4" resultid="1880"/><RANKING place="3" resultid="1881"/><RANKING place="5" resultid="1883"/><RANKING place="6" resultid="1888"/><RANKING place="2" resultid="1903"/><RANKING place="1" resultid="1922"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="270002" agemax="9" agemin="9" gender="F" name="Jahrgang 2016"><RANKINGS><RANKING place="11" resultid="1869"/><RANKING place="12" resultid="1870"/><RANKING place="9" resultid="1871"/><RANKING place="10" resultid="1878"/><RANKING place="13" resultid="1882"/><RANKING place="8" resultid="1891"/><RANKING place="4" resultid="1897"/><RANKING place="5" resultid="1902"/><RANKING place="7" resultid="1906"/><RANKING place="6" resultid="1910"/><RANKING place="2" resultid="1916"/><RANKING place="1" resultid="1923"/><RANKING place="3" resultid="1930"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="270003" agemax="10" agemin="10" gender="F" name="Jahrgang 2015"><RANKINGS><RANKING place="21" resultid="1864"/><RANKING place="20" resultid="1866"/><RANKING place="5" resultid="1873"/><RANKING place="16" resultid="1879"/><RANKING place="17" resultid="1884"/><RANKING place="12" resultid="1886"/><RANKING place="13" resultid="1889"/><RANKING place="18" resultid="1892"/><RANKING place="15" resultid="1893"/><RANKING place="7" resultid="1898"/><RANKING place="19" resultid="1899"/><RANKING place="-1" resultid="1900"/><RANKING place="9" resultid="1904"/><RANKING place="7" resultid="1909"/><RANKING place="10" resultid="1913"/><RANKING place="14" resultid="1915"/><RANKING place="11" resultid="1918"/><RANKING place="3" resultid="1925"/><RANKING place="4" resultid="1927"/><RANKING place="6" resultid="1929"/><RANKING place="-1" resultid="1931"/><RANKING place="1" resultid="1935"/><RANKING place="2" resultid="1947"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="270004" agemax="11" agemin="11" gender="F" name="Jahrgang 2014"><RANKINGS><RANKING place="15" resultid="1863"/><RANKING place="10" resultid="1865"/><RANKING place="13" resultid="1885"/><RANKING place="14" resultid="1887"/><RANKING place="12" resultid="1890"/><RANKING place="9" resultid="1905"/><RANKING place="11" resultid="1907"/><RANKING place="7" resultid="1908"/><RANKING place="5" resultid="1917"/><RANKING place="8" resultid="1919"/><RANKING place="6" resultid="1928"/><RANKING place="4" resultid="1936"/><RANKING place="2" resultid="1937"/><RANKING place="3" resultid="1963"/><RANKING place="1" resultid="1980"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="270005" agemax="12" agemin="12" gender="F" name="Jahrgang 2013"><RANKINGS><RANKING place="18" resultid="1862"/><RANKING place="-1" resultid="1872"/><RANKING place="-1" resultid="1875"/><RANKING place="16" resultid="1876"/><RANKING place="17" resultid="1877"/><RANKING place="13" resultid="1894"/><RANKING place="12" resultid="1896"/><RANKING place="14" resultid="1901"/><RANKING place="15" resultid="1912"/><RANKING place="-1" resultid="1914"/><RANKING place="11" resultid="1921"/><RANKING place="10" resultid="1924"/><RANKING place="8" resultid="1926"/><RANKING place="9" resultid="1933"/><RANKING place="7" resultid="1934"/><RANKING place="6" resultid="1938"/><RANKING place="5" resultid="1942"/><RANKING place="4" resultid="1960"/><RANKING place="1" resultid="1971"/><RANKING place="3" resultid="1982"/><RANKING place="2" resultid="1988"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="270006" agemax="13" agemin="13" gender="F" name="Jahrgang 2012"><RANKINGS><RANKING place="14" resultid="1867"/><RANKING place="11" resultid="1911"/><RANKING place="13" resultid="1939"/><RANKING place="12" resultid="1941"/><RANKING place="10" resultid="1944"/><RANKING place="7" resultid="1950"/><RANKING place="9" resultid="1951"/><RANKING place="4" resultid="1957"/><RANKING place="3" resultid="1959"/><RANKING place="8" resultid="1961"/><RANKING place="1" resultid="1969"/><RANKING place="2" resultid="1973"/><RANKING place="5" resultid="1986"/><RANKING place="6" resultid="1995"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="270007" agemax="14" agemin="14" gender="F" name="Jahrgang 2011"><RANKINGS><RANKING place="19" resultid="1895"/><RANKING place="18" resultid="1920"/><RANKING place="10" resultid="1945"/><RANKING place="13" resultid="1946"/><RANKING place="17" resultid="1948"/><RANKING place="14" resultid="1949"/><RANKING place="12" resultid="1953"/><RANKING place="20" resultid="1955"/><RANKING place="15" resultid="1962"/><RANKING place="-1" resultid="1970"/><RANKING place="7" resultid="1972"/><RANKING place="11" resultid="1981"/><RANKING place="16" resultid="1987"/><RANKING place="5" resultid="1990"/><RANKING place="8" resultid="1996"/><RANKING place="9" resultid="2000"/><RANKING place="6" resultid="2001"/><RANKING place="2" resultid="2004"/><RANKING place="3" resultid="2005"/><RANKING place="4" resultid="2016"/><RANKING place="1" resultid="2020"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="270008" agemax="15" agemin="15" gender="F" name="Jahrgang 2010"><RANKINGS><RANKING place="14" resultid="1940"/><RANKING place="15" resultid="1954"/><RANKING place="12" resultid="1964"/><RANKING place="10" resultid="1968"/><RANKING place="9" resultid="1976"/><RANKING place="13" resultid="1977"/><RANKING place="11" resultid="1978"/><RANKING place="6" resultid="1983"/><RANKING place="-1" resultid="1984"/><RANKING place="7" resultid="1985"/><RANKING place="4" resultid="1993"/><RANKING place="8" resultid="2002"/><RANKING place="3" resultid="2003"/><RANKING place="2" resultid="2007"/><RANKING place="5" resultid="2015"/><RANKING place="1" resultid="2018"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="270009" agemax="16" agemin="16" gender="F" name="Jahrgang 2009"><RANKINGS><RANKING place="-1" resultid="1932"/><RANKING place="15" resultid="1943"/><RANKING place="12" resultid="1952"/><RANKING place="16" resultid="1956"/><RANKING place="11" resultid="1958"/><RANKING place="14" resultid="1965"/><RANKING place="8" resultid="1966"/><RANKING place="13" resultid="1974"/><RANKING place="-1" resultid="1975"/><RANKING place="9" resultid="1992"/><RANKING place="10" resultid="1994"/><RANKING place="6" resultid="1997"/><RANKING place="7" resultid="1998"/><RANKING place="3" resultid="2006"/><RANKING place="5" resultid="2011"/><RANKING place="-1" resultid="2013"/><RANKING place="1" resultid="2021"/><RANKING place="2" resultid="2023"/><RANKING place="4" resultid="2024"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="270010" agemax="17" agemin="17" gender="F" name="Jahrgang 2008"><RANKINGS><RANKING place="3" resultid="1979"/><RANKING place="1" resultid="1989"/><RANKING place="-1" resultid="2009"/><RANKING place="2" resultid="2010"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="270011" agemax="-1" agemin="18" gender="F" name="Jahrgang 2007 und älter"><RANKINGS><RANKING place="8" resultid="1967"/><RANKING place="7" resultid="1991"/><RANKING place="5" resultid="1999"/><RANKING place="4" resultid="2008"/><RANKING place="-1" resultid="2012"/><RANKING place="3" resultid="2014"/><RANKING place="6" resultid="2017"/><RANKING place="2" resultid="2019"/><RANKING place="1" resultid="2022"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="252" number="1" order="1" status="OFFICIAL"/><HEAT heatid="253" number="2" order="2" status="OFFICIAL"/><HEAT heatid="254" number="3" order="3" status="OFFICIAL"/><HEAT heatid="255" number="4" order="4" status="OFFICIAL"/><HEAT heatid="256" number="5" order="5" status="OFFICIAL"/><HEAT heatid="257" number="6" order="6" status="OFFICIAL"/><HEAT heatid="258" number="7" order="7" status="OFFICIAL"/><HEAT heatid="259" number="8" order="8" status="OFFICIAL"/><HEAT heatid="260" number="9" order="9" status="OFFICIAL"/><HEAT heatid="261" number="10" order="10" status="OFFICIAL"/><HEAT heatid="262" number="11" order="11" status="OFFICIAL"/><HEAT heatid="263" number="12" order="12" status="OFFICIAL"/><HEAT heatid="264" number="13" order="13" status="OFFICIAL"/><HEAT heatid="265" number="14" order="14" status="OFFICIAL"/><HEAT heatid="266" number="15" order="15" status="OFFICIAL"/><HEAT heatid="267" number="16" order="16" status="OFFICIAL"/><HEAT heatid="268" number="17" order="17" status="OFFICIAL"/><HEAT heatid="269" number="18" order="18" status="OFFICIAL"/><HEAT heatid="270" number="19" order="19" status="OFFICIAL"/><HEAT heatid="271" number="20" order="20" status="OFFICIAL"/><HEAT heatid="272" number="21" order="21" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT><EVENT eventid="28" gender="M" number="28" order="28" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="700"/><SWIMSTYLE distance="50" name="50m Rücken Männer" relaycount="1" stroke="BACK"/><AGEGROUPS><AGEGROUP agegroupid="280001" agemax="8" agemin="8" gender="M" name="Jahrgang 2017"><RANKINGS><RANKING place="1" resultid="2037"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="280002" agemax="9" agemin="9" gender="M" name="Jahrgang 2016"><RANKINGS><RANKING place="9" resultid="2027"/><RANKING place="7" resultid="2031"/><RANKING place="6" resultid="2032"/><RANKING place="4" resultid="2033"/><RANKING place="3" resultid="2035"/><RANKING place="8" resultid="2038"/><RANKING place="5" resultid="2039"/><RANKING place="1" resultid="2053"/><RANKING place="2" resultid="2060"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="280003" agemax="10" agemin="10" gender="M" name="Jahrgang 2015"><RANKINGS><RANKING place="-1" resultid="2026"/><RANKING place="7" resultid="2034"/><RANKING place="12" resultid="2036"/><RANKING place="9" resultid="2040"/><RANKING place="6" resultid="2042"/><RANKING place="5" resultid="2044"/><RANKING place="13" resultid="2050"/><RANKING place="3" resultid="2058"/><RANKING place="10" resultid="2059"/><RANKING place="11" resultid="2061"/><RANKING place="8" resultid="2068"/><RANKING place="2" resultid="2069"/><RANKING place="1" resultid="2072"/><RANKING place="4" resultid="2084"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="280004" agemax="11" agemin="11" gender="M" name="Jahrgang 2014"><RANKINGS><RANKING place="12" resultid="2041"/><RANKING place="15" resultid="2046"/><RANKING place="14" resultid="2048"/><RANKING place="10" resultid="2051"/><RANKING place="5" resultid="2052"/><RANKING place="7" resultid="2055"/><RANKING place="13" resultid="2056"/><RANKING place="11" resultid="2057"/><RANKING place="6" resultid="2063"/><RANKING place="9" resultid="2065"/><RANKING place="4" resultid="2066"/><RANKING place="8" resultid="2067"/><RANKING place="2" resultid="2073"/><RANKING place="3" resultid="2074"/><RANKING place="1" resultid="2083"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="280005" agemax="12" agemin="12" gender="M" name="Jahrgang 2013"><RANKINGS><RANKING place="9" resultid="2029"/><RANKING place="-1" resultid="2043"/><RANKING place="7" resultid="2047"/><RANKING place="8" resultid="2049"/><RANKING place="6" resultid="2062"/><RANKING place="3" resultid="2075"/><RANKING place="4" resultid="2078"/><RANKING place="5" resultid="2087"/><RANKING place="1" resultid="2089"/><RANKING place="2" resultid="2092"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="280006" agemax="13" agemin="13" gender="M" name="Jahrgang 2012"><RANKINGS><RANKING place="9" resultid="2030"/><RANKING place="10" resultid="2054"/><RANKING place="8" resultid="2070"/><RANKING place="7" resultid="2071"/><RANKING place="-1" resultid="2076"/><RANKING place="5" resultid="2077"/><RANKING place="3" resultid="2079"/><RANKING place="6" resultid="2088"/><RANKING place="2" resultid="2096"/><RANKING place="1" resultid="2099"/><RANKING place="4" resultid="2101"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="280007" agemax="14" agemin="14" gender="M" name="Jahrgang 2011"><RANKINGS><RANKING place="17" resultid="2028"/><RANKING place="16" resultid="2045"/><RANKING place="15" resultid="2064"/><RANKING place="10" resultid="2080"/><RANKING place="5" resultid="2081"/><RANKING place="12" resultid="2085"/><RANKING place="13" resultid="2086"/><RANKING place="-1" resultid="2090"/><RANKING place="9" resultid="2091"/><RANKING place="11" resultid="2094"/><RANKING place="8" resultid="2095"/><RANKING place="-1" resultid="2097"/><RANKING place="4" resultid="2098"/><RANKING place="14" resultid="2100"/><RANKING place="2" resultid="2103"/><RANKING place="7" resultid="2106"/><RANKING place="6" resultid="2107"/><RANKING place="1" resultid="2110"/><RANKING place="3" resultid="2113"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="280008" agemax="15" agemin="15" gender="M" name="Jahrgang 2010"><RANKINGS><RANKING place="11" resultid="2025"/><RANKING place="-1" resultid="2082"/><RANKING place="8" resultid="2093"/><RANKING place="9" resultid="2102"/><RANKING place="6" resultid="2105"/><RANKING place="10" resultid="2108"/><RANKING place="7" resultid="2109"/><RANKING place="-1" resultid="2114"/><RANKING place="5" resultid="2116"/><RANKING place="4" resultid="2121"/><RANKING place="3" resultid="2125"/><RANKING place="1" resultid="2128"/><RANKING place="2" resultid="2137"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="280009" agemax="16" agemin="16" gender="M" name="Jahrgang 2009"><RANKINGS><RANKING place="9" resultid="2104"/><RANKING place="7" resultid="2111"/><RANKING place="6" resultid="2112"/><RANKING place="8" resultid="2115"/><RANKING place="-1" resultid="2117"/><RANKING place="4" resultid="2119"/><RANKING place="5" resultid="2122"/><RANKING place="-1" resultid="2124"/><RANKING place="2" resultid="2127"/><RANKING place="3" resultid="2132"/><RANKING place="1" resultid="2136"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="280010" agemax="17" agemin="17" gender="M" name="Jahrgang 2008"><RANKINGS><RANKING place="-1" resultid="2129"/><RANKING place="2" resultid="2130"/><RANKING place="1" resultid="2135"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="280011" agemax="-1" agemin="18" gender="M" name="Jahrgang 2007 und älter"><RANKINGS><RANKING place="-1" resultid="2118"/><RANKING place="4" resultid="2120"/><RANKING place="5" resultid="2123"/><RANKING place="3" resultid="2126"/><RANKING place="6" resultid="2131"/><RANKING place="1" resultid="2133"/><RANKING place="2" resultid="2134"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="273" number="1" order="1" status="OFFICIAL"/><HEAT heatid="274" number="2" order="2" status="OFFICIAL"/><HEAT heatid="275" number="3" order="3" status="OFFICIAL"/><HEAT heatid="276" number="4" order="4" status="OFFICIAL"/><HEAT heatid="277" number="5" order="5" status="OFFICIAL"/><HEAT heatid="278" number="6" order="6" status="OFFICIAL"/><HEAT heatid="279" number="7" order="7" status="OFFICIAL"/><HEAT heatid="280" number="8" order="8" status="OFFICIAL"/><HEAT heatid="281" number="9" order="9" status="OFFICIAL"/><HEAT heatid="282" number="10" order="10" status="OFFICIAL"/><HEAT heatid="283" number="11" order="11" status="OFFICIAL"/><HEAT heatid="284" number="12" order="12" status="OFFICIAL"/><HEAT heatid="285" number="13" order="13" status="OFFICIAL"/><HEAT heatid="286" number="14" order="14" status="OFFICIAL"/><HEAT heatid="287" number="15" order="15" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT><EVENT eventid="29" gender="F" number="29" order="29" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="700"/><SWIMSTYLE distance="200" name="200m Freistil Frauen" relaycount="1" stroke="FREE"/><AGEGROUPS><AGEGROUP agegroupid="290001" agemax="9" agemin="9" gender="F" name="Jahrgang 2016"><RANKINGS><RANKING place="6" resultid="2141"/><RANKING place="8" resultid="2152"/><RANKING place="5" resultid="2155"/><RANKING place="7" resultid="2157"/><RANKING place="3" resultid="2166"/><RANKING place="1" resultid="2178"/><RANKING place="4" resultid="2179"/><RANKING place="2" resultid="2181"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="290002" agemax="10" agemin="10" gender="F" name="Jahrgang 2015"><RANKINGS><RANKING place="11" resultid="2139"/><RANKING place="12" resultid="2140"/><RANKING place="-1" resultid="2142"/><RANKING place="9" resultid="2146"/><RANKING place="10" resultid="2150"/><RANKING place="2" resultid="2154"/><RANKING place="8" resultid="2161"/><RANKING place="7" resultid="2163"/><RANKING place="6" resultid="2165"/><RANKING place="4" resultid="2176"/><RANKING place="5" resultid="2182"/><RANKING place="1" resultid="2203"/><RANKING place="3" resultid="2213"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="290003" agemax="11" agemin="11" gender="F" name="Jahrgang 2014"><RANKINGS><RANKING place="27" resultid="2138"/><RANKING place="23" resultid="2144"/><RANKING place="20" resultid="2147"/><RANKING place="25" resultid="2148"/><RANKING place="28" resultid="2149"/><RANKING place="21" resultid="2151"/><RANKING place="26" resultid="2156"/><RANKING place="24" resultid="2158"/><RANKING place="15" resultid="2160"/><RANKING place="19" resultid="2162"/><RANKING place="22" resultid="2167"/><RANKING place="9" resultid="2169"/><RANKING place="17" resultid="2171"/><RANKING place="16" resultid="2174"/><RANKING place="12" resultid="2175"/><RANKING place="18" resultid="2177"/><RANKING place="10" resultid="2184"/><RANKING place="11" resultid="2186"/><RANKING place="13" resultid="2188"/><RANKING place="14" resultid="2189"/><RANKING place="5" resultid="2194"/><RANKING place="4" resultid="2204"/><RANKING place="3" resultid="2209"/><RANKING place="6" resultid="2210"/><RANKING place="2" resultid="2211"/><RANKING place="7" resultid="2212"/><RANKING place="1" resultid="2220"/><RANKING place="8" resultid="2229"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="290004" agemax="12" agemin="12" gender="F" name="Jahrgang 2013"><RANKINGS><RANKING place="18" resultid="2143"/><RANKING place="-1" resultid="2145"/><RANKING place="13" resultid="2153"/><RANKING place="17" resultid="2159"/><RANKING place="16" resultid="2164"/><RANKING place="15" resultid="2168"/><RANKING place="14" resultid="2170"/><RANKING place="11" resultid="2187"/><RANKING place="10" resultid="2190"/><RANKING place="9" resultid="2191"/><RANKING place="12" resultid="2196"/><RANKING place="8" resultid="2199"/><RANKING place="4" resultid="2200"/><RANKING place="7" resultid="2202"/><RANKING place="6" resultid="2215"/><RANKING place="-1" resultid="2219"/><RANKING place="3" resultid="2223"/><RANKING place="2" resultid="2233"/><RANKING place="5" resultid="2241"/><RANKING place="1" resultid="2252"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="290005" agemax="13" agemin="13" gender="F" name="Jahrgang 2012"><RANKINGS><RANKING place="14" resultid="2185"/><RANKING place="13" resultid="2195"/><RANKING place="12" resultid="2206"/><RANKING place="11" resultid="2216"/><RANKING place="10" resultid="2217"/><RANKING place="9" resultid="2221"/><RANKING place="7" resultid="2232"/><RANKING place="8" resultid="2237"/><RANKING place="6" resultid="2240"/><RANKING place="3" resultid="2243"/><RANKING place="4" resultid="2249"/><RANKING place="5" resultid="2250"/><RANKING place="2" resultid="2256"/><RANKING place="1" resultid="2282"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="290006" agemax="14" agemin="14" gender="F" name="Jahrgang 2011"><RANKINGS><RANKING place="17" resultid="2173"/><RANKING place="19" resultid="2192"/><RANKING place="16" resultid="2193"/><RANKING place="15" resultid="2198"/><RANKING place="14" resultid="2214"/><RANKING place="18" resultid="2224"/><RANKING place="13" resultid="2225"/><RANKING place="6" resultid="2239"/><RANKING place="10" resultid="2242"/><RANKING place="12" resultid="2245"/><RANKING place="11" resultid="2248"/><RANKING place="8" resultid="2258"/><RANKING place="7" resultid="2262"/><RANKING place="5" resultid="2266"/><RANKING place="9" resultid="2267"/><RANKING place="4" resultid="2270"/><RANKING place="3" resultid="2274"/><RANKING place="2" resultid="2276"/><RANKING place="1" resultid="2281"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="290007" agemax="15" agemin="15" gender="F" name="Jahrgang 2010"><RANKINGS><RANKING place="14" resultid="2172"/><RANKING place="11" resultid="2218"/><RANKING place="-1" resultid="2222"/><RANKING place="9" resultid="2227"/><RANKING place="12" resultid="2228"/><RANKING place="7" resultid="2231"/><RANKING place="10" resultid="2236"/><RANKING place="6" resultid="2244"/><RANKING place="13" resultid="2251"/><RANKING place="3" resultid="2253"/><RANKING place="8" resultid="2259"/><RANKING place="5" resultid="2269"/><RANKING place="2" resultid="2273"/><RANKING place="4" resultid="2279"/><RANKING place="1" resultid="2287"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="290008" agemax="16" agemin="16" gender="F" name="Jahrgang 2009"><RANKINGS><RANKING place="12" resultid="2183"/><RANKING place="-1" resultid="2197"/><RANKING place="14" resultid="2201"/><RANKING place="16" resultid="2205"/><RANKING place="13" resultid="2208"/><RANKING place="15" resultid="2230"/><RANKING place="11" resultid="2234"/><RANKING place="8" resultid="2246"/><RANKING place="10" resultid="2247"/><RANKING place="6" resultid="2254"/><RANKING place="7" resultid="2255"/><RANKING place="5" resultid="2257"/><RANKING place="9" resultid="2260"/><RANKING place="3" resultid="2264"/><RANKING place="4" resultid="2268"/><RANKING place="-1" resultid="2277"/><RANKING place="2" resultid="2278"/><RANKING place="1" resultid="2289"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="290009" agemax="17" agemin="17" gender="F" name="Jahrgang 2008"><RANKINGS><RANKING place="7" resultid="2235"/><RANKING place="6" resultid="2261"/><RANKING place="4" resultid="2263"/><RANKING place="5" resultid="2275"/><RANKING place="3" resultid="2283"/><RANKING place="1" resultid="2284"/><RANKING place="2" resultid="2290"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="290010" agemax="-1" agemin="18" gender="F" name="Jahrgang 2007 und älter"><RANKINGS><RANKING place="11" resultid="2180"/><RANKING place="10" resultid="2207"/><RANKING place="9" resultid="2226"/><RANKING place="7" resultid="2238"/><RANKING place="8" resultid="2265"/><RANKING place="4" resultid="2271"/><RANKING place="5" resultid="2272"/><RANKING place="6" resultid="2280"/><RANKING place="3" resultid="2285"/><RANKING place="2" resultid="2286"/><RANKING place="1" resultid="2288"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="288" number="1" order="1" status="OFFICIAL"/><HEAT heatid="289" number="2" order="2" status="OFFICIAL"/><HEAT heatid="290" number="3" order="3" status="OFFICIAL"/><HEAT heatid="291" number="4" order="4" status="OFFICIAL"/><HEAT heatid="292" number="5" order="5" status="OFFICIAL"/><HEAT heatid="293" number="6" order="6" status="OFFICIAL"/><HEAT heatid="294" number="7" order="7" status="OFFICIAL"/><HEAT heatid="295" number="8" order="8" status="OFFICIAL"/><HEAT heatid="296" number="9" order="9" status="OFFICIAL"/><HEAT heatid="297" number="10" order="10" status="OFFICIAL"/><HEAT heatid="298" number="11" order="11" status="OFFICIAL"/><HEAT heatid="299" number="12" order="12" status="OFFICIAL"/><HEAT heatid="300" number="13" order="13" status="OFFICIAL"/><HEAT heatid="301" number="14" order="14" status="OFFICIAL"/><HEAT heatid="302" number="15" order="15" status="OFFICIAL"/><HEAT heatid="303" number="16" order="16" status="OFFICIAL"/><HEAT heatid="304" number="17" order="17" status="OFFICIAL"/><HEAT heatid="305" number="18" order="18" status="OFFICIAL"/><HEAT heatid="306" number="19" order="19" status="OFFICIAL"/><HEAT heatid="307" number="20" order="20" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT><EVENT eventid="30" gender="M" number="30" order="30" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="700"/><SWIMSTYLE distance="200" name="200m Freistil Männer" relaycount="1" stroke="FREE"/><AGEGROUPS><AGEGROUP agegroupid="300001" agemax="9" agemin="9" gender="M" name="Jahrgang 2016"><RANKINGS><RANKING place="4" resultid="2297"/><RANKING place="5" resultid="2298"/><RANKING place="3" resultid="2300"/><RANKING place="2" resultid="2308"/><RANKING place="1" resultid="2333"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="300002" agemax="10" agemin="10" gender="M" name="Jahrgang 2015"><RANKINGS><RANKING place="16" resultid="2291"/><RANKING place="-1" resultid="2294"/><RANKING place="18" resultid="2301"/><RANKING place="19" resultid="2302"/><RANKING place="13" resultid="2304"/><RANKING place="15" resultid="2306"/><RANKING place="17" resultid="2311"/><RANKING place="11" resultid="2316"/><RANKING place="14" resultid="2317"/><RANKING place="12" resultid="2318"/><RANKING place="2" resultid="2322"/><RANKING place="6" resultid="2323"/><RANKING place="10" resultid="2325"/><RANKING place="4" resultid="2326"/><RANKING place="8" resultid="2328"/><RANKING place="9" resultid="2329"/><RANKING place="7" resultid="2332"/><RANKING place="3" resultid="2334"/><RANKING place="1" resultid="2338"/><RANKING place="5" resultid="2346"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="300003" agemax="11" agemin="11" gender="M" name="Jahrgang 2014"><RANKINGS><RANKING place="15" resultid="2299"/><RANKING place="14" resultid="2303"/><RANKING place="13" resultid="2305"/><RANKING place="11" resultid="2314"/><RANKING place="10" resultid="2315"/><RANKING place="9" resultid="2319"/><RANKING place="6" resultid="2320"/><RANKING place="8" resultid="2327"/><RANKING place="5" resultid="2336"/><RANKING place="7" resultid="2340"/><RANKING place="12" resultid="2342"/><RANKING place="4" resultid="2350"/><RANKING place="3" resultid="2353"/><RANKING place="2" resultid="2358"/><RANKING place="1" resultid="2362"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="300004" agemax="12" agemin="12" gender="M" name="Jahrgang 2013"><RANKINGS><RANKING place="18" resultid="2296"/><RANKING place="16" resultid="2307"/><RANKING place="-1" resultid="2309"/><RANKING place="19" resultid="2310"/><RANKING place="17" resultid="2312"/><RANKING place="14" resultid="2331"/><RANKING place="13" resultid="2335"/><RANKING place="12" resultid="2337"/><RANKING place="15" resultid="2339"/><RANKING place="10" resultid="2341"/><RANKING place="6" resultid="2343"/><RANKING place="11" resultid="2344"/><RANKING place="9" resultid="2345"/><RANKING place="8" resultid="2351"/><RANKING place="2" resultid="2355"/><RANKING place="4" resultid="2360"/><RANKING place="7" resultid="2365"/><RANKING place="5" resultid="2367"/><RANKING place="3" resultid="2378"/><RANKING place="1" resultid="2388"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="300005" agemax="13" agemin="13" gender="M" name="Jahrgang 2012"><RANKINGS><RANKING place="10" resultid="2295"/><RANKING place="8" resultid="2321"/><RANKING place="9" resultid="2349"/><RANKING place="4" resultid="2352"/><RANKING place="7" resultid="2372"/><RANKING place="6" resultid="2374"/><RANKING place="5" resultid="2377"/><RANKING place="2" resultid="2381"/><RANKING place="3" resultid="2386"/><RANKING place="1" resultid="2402"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="300006" agemax="14" agemin="14" gender="M" name="Jahrgang 2011"><RANKINGS><RANKING place="23" resultid="2292"/><RANKING place="22" resultid="2313"/><RANKING place="21" resultid="2324"/><RANKING place="20" resultid="2330"/><RANKING place="19" resultid="2348"/><RANKING place="18" resultid="2354"/><RANKING place="17" resultid="2356"/><RANKING place="-1" resultid="2357"/><RANKING place="16" resultid="2361"/><RANKING place="13" resultid="2363"/><RANKING place="11" resultid="2368"/><RANKING place="15" resultid="2370"/><RANKING place="14" resultid="2373"/><RANKING place="8" resultid="2380"/><RANKING place="9" resultid="2382"/><RANKING place="-1" resultid="2383"/><RANKING place="7" resultid="2387"/><RANKING place="5" resultid="2393"/><RANKING place="6" resultid="2394"/><RANKING place="12" resultid="2395"/><RANKING place="4" resultid="2396"/><RANKING place="2" resultid="2400"/><RANKING place="10" resultid="2403"/><RANKING place="3" resultid="2404"/><RANKING place="1" resultid="2408"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="300007" agemax="15" agemin="15" gender="M" name="Jahrgang 2010"><RANKINGS><RANKING place="15" resultid="2293"/><RANKING place="16" resultid="2347"/><RANKING place="11" resultid="2364"/><RANKING place="14" resultid="2366"/><RANKING place="-1" resultid="2375"/><RANKING place="12" resultid="2379"/><RANKING place="10" resultid="2384"/><RANKING place="13" resultid="2389"/><RANKING place="9" resultid="2391"/><RANKING place="8" resultid="2392"/><RANKING place="5" resultid="2398"/><RANKING place="7" resultid="2399"/><RANKING place="6" resultid="2405"/><RANKING place="2" resultid="2406"/><RANKING place="4" resultid="2407"/><RANKING place="3" resultid="2411"/><RANKING place="1" resultid="2422"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="300008" agemax="16" agemin="16" gender="M" name="Jahrgang 2009"><RANKINGS><RANKING place="13" resultid="2369"/><RANKING place="12" resultid="2371"/><RANKING place="10" resultid="2376"/><RANKING place="11" resultid="2385"/><RANKING place="9" resultid="2390"/><RANKING place="8" resultid="2401"/><RANKING place="5" resultid="2409"/><RANKING place="2" resultid="2413"/><RANKING place="7" resultid="2415"/><RANKING place="3" resultid="2416"/><RANKING place="4" resultid="2418"/><RANKING place="1" resultid="2419"/><RANKING place="6" resultid="2425"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="300009" agemax="17" agemin="17" gender="M" name="Jahrgang 2008"><RANKINGS><RANKING place="2" resultid="2359"/><RANKING place="-1" resultid="2410"/><RANKING place="1" resultid="2412"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="300010" agemax="-1" agemin="18" gender="M" name="Jahrgang 2007 und älter"><RANKINGS><RANKING place="6" resultid="2397"/><RANKING place="4" resultid="2414"/><RANKING place="3" resultid="2417"/><RANKING place="2" resultid="2420"/><RANKING place="1" resultid="2421"/><RANKING place="5" resultid="2423"/><RANKING place="7" resultid="2424"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="308" number="1" order="1" status="OFFICIAL"/><HEAT heatid="309" number="2" order="2" status="OFFICIAL"/><HEAT heatid="310" number="3" order="3" status="OFFICIAL"/><HEAT heatid="311" number="4" order="4" status="OFFICIAL"/><HEAT heatid="312" number="5" order="5" status="OFFICIAL"/><HEAT heatid="313" number="6" order="6" status="OFFICIAL"/><HEAT heatid="314" number="7" order="7" status="OFFICIAL"/><HEAT heatid="315" number="8" order="8" status="OFFICIAL"/><HEAT heatid="316" number="9" order="9" status="OFFICIAL"/><HEAT heatid="317" number="10" order="10" status="OFFICIAL"/><HEAT heatid="318" number="11" order="11" status="OFFICIAL"/><HEAT heatid="319" number="12" order="12" status="OFFICIAL"/><HEAT heatid="320" number="13" order="13" status="OFFICIAL"/><HEAT heatid="321" number="14" order="14" status="OFFICIAL"/><HEAT heatid="322" number="15" order="15" status="OFFICIAL"/><HEAT heatid="323" number="16" order="16" status="OFFICIAL"/><HEAT heatid="324" number="17" order="17" status="OFFICIAL"/><HEAT heatid="325" number="18" order="18" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT><EVENT eventid="31" gender="F" number="31" order="31" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="700"/><SWIMSTYLE distance="100" name="100m Brust Frauen" relaycount="1" stroke="BREAST"/><AGEGROUPS><AGEGROUP agegroupid="310001" agemax="9" agemin="9" gender="F" name="Jahrgang 2016"><RANKINGS><RANKING place="6" resultid="2436"/><RANKING place="5" resultid="2438"/><RANKING place="8" resultid="2440"/><RANKING place="7" resultid="2443"/><RANKING place="4" resultid="2454"/><RANKING place="2" resultid="2461"/><RANKING place="3" resultid="2465"/><RANKING place="1" resultid="2474"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="310002" agemax="10" agemin="10" gender="F" name="Jahrgang 2015"><RANKINGS><RANKING place="18" resultid="2428"/><RANKING place="13" resultid="2431"/><RANKING place="17" resultid="2433"/><RANKING place="15" resultid="2444"/><RANKING place="-1" resultid="2445"/><RANKING place="4" resultid="2446"/><RANKING place="12" resultid="2447"/><RANKING place="16" resultid="2452"/><RANKING place="11" resultid="2455"/><RANKING place="14" resultid="2458"/><RANKING place="-1" resultid="2459"/><RANKING place="6" resultid="2460"/><RANKING place="10" resultid="2462"/><RANKING place="8" resultid="2467"/><RANKING place="9" resultid="2468"/><RANKING place="7" resultid="2471"/><RANKING place="5" resultid="2480"/><RANKING place="3" resultid="2482"/><RANKING place="2" resultid="2484"/><RANKING place="1" resultid="2494"/><RANKING place="-1" resultid="2511"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="310003" agemax="11" agemin="11" gender="F" name="Jahrgang 2014"><RANKINGS><RANKING place="24" resultid="2427"/><RANKING place="22" resultid="2435"/><RANKING place="23" resultid="2439"/><RANKING place="18" resultid="2441"/><RANKING place="20" resultid="2442"/><RANKING place="19" resultid="2448"/><RANKING place="21" resultid="2449"/><RANKING place="17" resultid="2451"/><RANKING place="15" resultid="2464"/><RANKING place="13" resultid="2469"/><RANKING place="12" resultid="2470"/><RANKING place="10" resultid="2476"/><RANKING place="14" resultid="2477"/><RANKING place="16" resultid="2478"/><RANKING place="6" resultid="2481"/><RANKING place="-1" resultid="2485"/><RANKING place="9" resultid="2486"/><RANKING place="4" resultid="2487"/><RANKING place="11" resultid="2489"/><RANKING place="7" resultid="2491"/><RANKING place="5" resultid="2492"/><RANKING place="8" resultid="2497"/><RANKING place="2" resultid="2498"/><RANKING place="3" resultid="2506"/><RANKING place="1" resultid="2512"/><RANKING place="-1" resultid="2522"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="310004" agemax="12" agemin="12" gender="F" name="Jahrgang 2013"><RANKINGS><RANKING place="26" resultid="2426"/><RANKING place="25" resultid="2429"/><RANKING place="-1" resultid="2430"/><RANKING place="27" resultid="2432"/><RANKING place="21" resultid="2437"/><RANKING place="24" resultid="2450"/><RANKING place="16" resultid="2453"/><RANKING place="20" resultid="2456"/><RANKING place="-1" resultid="2457"/><RANKING place="11" resultid="2463"/><RANKING place="22" resultid="2466"/><RANKING place="23" resultid="2472"/><RANKING place="19" resultid="2473"/><RANKING place="18" resultid="2479"/><RANKING place="17" resultid="2483"/><RANKING place="-1" resultid="2488"/><RANKING place="12" resultid="2490"/><RANKING place="15" resultid="2496"/><RANKING place="-1" resultid="2499"/><RANKING place="14" resultid="2502"/><RANKING place="5" resultid="2503"/><RANKING place="10" resultid="2505"/><RANKING place="13" resultid="2507"/><RANKING place="8" resultid="2509"/><RANKING place="9" resultid="2517"/><RANKING place="4" resultid="2524"/><RANKING place="6" resultid="2530"/><RANKING place="3" resultid="2532"/><RANKING place="7" resultid="2533"/><RANKING place="2" resultid="2541"/><RANKING place="1" resultid="2544"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="310005" agemax="13" agemin="13" gender="F" name="Jahrgang 2012"><RANKINGS><RANKING place="11" resultid="2434"/><RANKING place="10" resultid="2500"/><RANKING place="9" resultid="2514"/><RANKING place="6" resultid="2518"/><RANKING place="8" resultid="2520"/><RANKING place="5" resultid="2526"/><RANKING place="7" resultid="2535"/><RANKING place="3" resultid="2539"/><RANKING place="4" resultid="2545"/><RANKING place="1" resultid="2556"/><RANKING place="2" resultid="2561"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="310006" agemax="14" agemin="14" gender="F" name="Jahrgang 2011"><RANKINGS><RANKING place="13" resultid="2495"/><RANKING place="12" resultid="2501"/><RANKING place="10" resultid="2508"/><RANKING place="11" resultid="2521"/><RANKING place="8" resultid="2525"/><RANKING place="9" resultid="2531"/><RANKING place="5" resultid="2534"/><RANKING place="6" resultid="2538"/><RANKING place="7" resultid="2546"/><RANKING place="2" resultid="2548"/><RANKING place="4" resultid="2550"/><RANKING place="3" resultid="2557"/><RANKING place="1" resultid="2564"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="310007" agemax="15" agemin="15" gender="F" name="Jahrgang 2010"><RANKINGS><RANKING place="9" resultid="2504"/><RANKING place="8" resultid="2510"/><RANKING place="7" resultid="2527"/><RANKING place="5" resultid="2528"/><RANKING place="6" resultid="2537"/><RANKING place="3" resultid="2553"/><RANKING place="4" resultid="2559"/><RANKING place="2" resultid="2560"/><RANKING place="1" resultid="2565"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="310008" agemax="16" agemin="16" gender="F" name="Jahrgang 2009"><RANKINGS><RANKING place="13" resultid="2475"/><RANKING place="12" resultid="2513"/><RANKING place="11" resultid="2515"/><RANKING place="-1" resultid="2519"/><RANKING place="10" resultid="2529"/><RANKING place="8" resultid="2549"/><RANKING place="6" resultid="2552"/><RANKING place="5" resultid="2555"/><RANKING place="4" resultid="2558"/><RANKING place="9" resultid="2562"/><RANKING place="2" resultid="2563"/><RANKING place="1" resultid="2566"/><RANKING place="7" resultid="2569"/><RANKING place="3" resultid="2570"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="310009" agemax="17" agemin="17" gender="F" name="Jahrgang 2008"><RANKINGS><RANKING place="1" resultid="2540"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="310010" agemax="-1" agemin="18" gender="F" name="Jahrgang 2007 und älter"><RANKINGS><RANKING place="11" resultid="2493"/><RANKING place="9" resultid="2516"/><RANKING place="10" resultid="2523"/><RANKING place="8" resultid="2536"/><RANKING place="3" resultid="2542"/><RANKING place="4" resultid="2543"/><RANKING place="5" resultid="2547"/><RANKING place="7" resultid="2551"/><RANKING place="6" resultid="2554"/><RANKING place="1" resultid="2567"/><RANKING place="2" resultid="2568"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="326" number="1" order="1" status="OFFICIAL"/><HEAT heatid="327" number="2" order="2" status="OFFICIAL"/><HEAT heatid="328" number="3" order="3" status="OFFICIAL"/><HEAT heatid="329" number="4" order="4" status="OFFICIAL"/><HEAT heatid="330" number="5" order="5" status="OFFICIAL"/><HEAT heatid="331" number="6" order="6" status="OFFICIAL"/><HEAT heatid="332" number="7" order="7" status="OFFICIAL"/><HEAT heatid="333" number="8" order="8" status="OFFICIAL"/><HEAT heatid="334" number="9" order="9" status="OFFICIAL"/><HEAT heatid="335" number="10" order="10" status="OFFICIAL"/><HEAT heatid="336" number="11" order="11" status="OFFICIAL"/><HEAT heatid="337" number="12" order="12" status="OFFICIAL"/><HEAT heatid="338" number="13" order="13" status="OFFICIAL"/><HEAT heatid="339" number="14" order="14" status="OFFICIAL"/><HEAT heatid="340" number="15" order="15" status="OFFICIAL"/><HEAT heatid="341" number="16" order="16" status="OFFICIAL"/><HEAT heatid="342" number="17" order="17" status="OFFICIAL"/><HEAT heatid="343" number="18" order="18" status="OFFICIAL"/><HEAT heatid="344" number="19" order="19" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT><EVENT eventid="32" gender="M" number="32" order="32" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="700"/><SWIMSTYLE distance="100" name="100m Brust Männer" relaycount="1" stroke="BREAST"/><AGEGROUPS><AGEGROUP agegroupid="320001" agemax="9" agemin="9" gender="M" name="Jahrgang 2016"><RANKINGS/></AGEGROUP><AGEGROUP agegroupid="320002" agemax="10" agemin="10" gender="M" name="Jahrgang 2015"><RANKINGS><RANKING place="8" resultid="2576"/><RANKING place="7" resultid="2579"/><RANKING place="11" resultid="2580"/><RANKING place="9" resultid="2582"/><RANKING place="10" resultid="2583"/><RANKING place="5" resultid="2590"/><RANKING place="6" resultid="2593"/><RANKING place="4" resultid="2598"/><RANKING place="2" resultid="2601"/><RANKING place="1" resultid="2602"/><RANKING place="3" resultid="2609"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="320003" agemax="11" agemin="11" gender="M" name="Jahrgang 2014"><RANKINGS><RANKING place="14" resultid="2577"/><RANKING place="15" resultid="2578"/><RANKING place="13" resultid="2581"/><RANKING place="10" resultid="2584"/><RANKING place="12" resultid="2586"/><RANKING place="11" resultid="2588"/><RANKING place="-1" resultid="2589"/><RANKING place="9" resultid="2591"/><RANKING place="4" resultid="2592"/><RANKING place="8" resultid="2594"/><RANKING place="6" resultid="2595"/><RANKING place="7" resultid="2596"/><RANKING place="5" resultid="2599"/><RANKING place="3" resultid="2600"/><RANKING place="2" resultid="2611"/><RANKING place="1" resultid="2612"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="320004" agemax="12" agemin="12" gender="M" name="Jahrgang 2013"><RANKINGS><RANKING place="7" resultid="2571"/><RANKING place="9" resultid="2573"/><RANKING place="8" resultid="2575"/><RANKING place="-1" resultid="2585"/><RANKING place="5" resultid="2587"/><RANKING place="4" resultid="2597"/><RANKING place="6" resultid="2604"/><RANKING place="3" resultid="2605"/><RANKING place="2" resultid="2607"/><RANKING place="1" resultid="2634"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="320005" agemax="13" agemin="13" gender="M" name="Jahrgang 2012"><RANKINGS><RANKING place="7" resultid="2574"/><RANKING place="6" resultid="2603"/><RANKING place="5" resultid="2606"/><RANKING place="3" resultid="2608"/><RANKING place="4" resultid="2610"/><RANKING place="2" resultid="2614"/><RANKING place="1" resultid="2627"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="320006" agemax="14" agemin="14" gender="M" name="Jahrgang 2011"><RANKINGS><RANKING place="15" resultid="2572"/><RANKING place="12" resultid="2613"/><RANKING place="11" resultid="2615"/><RANKING place="7" resultid="2616"/><RANKING place="14" resultid="2617"/><RANKING place="10" resultid="2618"/><RANKING place="13" resultid="2619"/><RANKING place="4" resultid="2620"/><RANKING place="6" resultid="2622"/><RANKING place="8" resultid="2623"/><RANKING place="5" resultid="2624"/><RANKING place="-1" resultid="2625"/><RANKING place="9" resultid="2626"/><RANKING place="3" resultid="2629"/><RANKING place="2" resultid="2632"/><RANKING place="-1" resultid="2637"/><RANKING place="1" resultid="2638"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="320007" agemax="15" agemin="15" gender="M" name="Jahrgang 2010"><RANKINGS><RANKING place="8" resultid="2621"/><RANKING place="7" resultid="2631"/><RANKING place="4" resultid="2633"/><RANKING place="3" resultid="2639"/><RANKING place="6" resultid="2642"/><RANKING place="5" resultid="2646"/><RANKING place="2" resultid="2648"/><RANKING place="1" resultid="2649"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="320008" agemax="16" agemin="16" gender="M" name="Jahrgang 2009"><RANKINGS><RANKING place="-1" resultid="2628"/><RANKING place="5" resultid="2630"/><RANKING place="2" resultid="2643"/><RANKING place="4" resultid="2650"/><RANKING place="3" resultid="2651"/><RANKING place="1" resultid="2654"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="320009" agemax="17" agemin="17" gender="M" name="Jahrgang 2008"><RANKINGS><RANKING place="5" resultid="2636"/><RANKING place="4" resultid="2640"/><RANKING place="3" resultid="2647"/><RANKING place="2" resultid="2652"/><RANKING place="1" resultid="2656"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="320010" agemax="-1" agemin="18" gender="M" name="Jahrgang 2007 und älter"><RANKINGS><RANKING place="7" resultid="2635"/><RANKING place="6" resultid="2641"/><RANKING place="1" resultid="2644"/><RANKING place="5" resultid="2645"/><RANKING place="3" resultid="2653"/><RANKING place="2" resultid="2655"/><RANKING place="4" resultid="2657"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="345" number="1" order="1" status="OFFICIAL"/><HEAT heatid="346" number="2" order="2" status="OFFICIAL"/><HEAT heatid="347" number="3" order="3" status="OFFICIAL"/><HEAT heatid="348" number="4" order="4" status="OFFICIAL"/><HEAT heatid="349" number="5" order="5" status="OFFICIAL"/><HEAT heatid="350" number="6" order="6" status="OFFICIAL"/><HEAT heatid="351" number="7" order="7" status="OFFICIAL"/><HEAT heatid="352" number="8" order="8" status="OFFICIAL"/><HEAT heatid="353" number="9" order="9" status="OFFICIAL"/><HEAT heatid="354" number="10" order="10" status="OFFICIAL"/><HEAT heatid="355" number="11" order="11" status="OFFICIAL"/><HEAT heatid="356" number="12" order="12" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT><EVENT eventid="33" gender="F" number="33" order="33" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="700"/><SWIMSTYLE distance="200" name="200m Schmetterling Frauen" relaycount="1" stroke="FLY"/><AGEGROUPS><AGEGROUP agegroupid="330001" agemax="11" agemin="11" gender="F" name="Jahrgang 2014"><RANKINGS><RANKING place="1" resultid="2666"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="330002" agemax="12" agemin="12" gender="F" name="Jahrgang 2013"><RANKINGS><RANKING place="3" resultid="2661"/><RANKING place="2" resultid="2662"/><RANKING place="1" resultid="2665"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="330003" agemax="13" agemin="13" gender="F" name="Jahrgang 2012"><RANKINGS><RANKING place="-1" resultid="2660"/><RANKING place="3" resultid="2664"/><RANKING place="1" resultid="2672"/><RANKING place="2" resultid="2674"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="330004" agemax="14" agemin="14" gender="F" name="Jahrgang 2011"><RANKINGS><RANKING place="4" resultid="2659"/><RANKING place="3" resultid="2663"/><RANKING place="2" resultid="2671"/><RANKING place="1" resultid="2676"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="330005" agemax="15" agemin="15" gender="F" name="Jahrgang 2010"><RANKINGS><RANKING place="2" resultid="2658"/><RANKING place="1" resultid="2682"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="330006" agemax="16" agemin="16" gender="F" name="Jahrgang 2009"><RANKINGS><RANKING place="-1" resultid="2667"/><RANKING place="2" resultid="2668"/><RANKING place="3" resultid="2670"/><RANKING place="1" resultid="2677"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="330007" agemax="17" agemin="17" gender="F" name="Jahrgang 2008"><RANKINGS><RANKING place="2" resultid="2679"/><RANKING place="1" resultid="2680"/><RANKING place="3" resultid="2681"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="330008" agemax="-1" agemin="18" gender="F" name="Jahrgang 2007 und älter"><RANKINGS><RANKING place="2" resultid="2669"/><RANKING place="4" resultid="2673"/><RANKING place="1" resultid="2675"/><RANKING place="3" resultid="2678"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="357" number="1" order="1" status="OFFICIAL"/><HEAT heatid="358" number="2" order="2" status="OFFICIAL"/><HEAT heatid="359" number="3" order="3" status="OFFICIAL"/><HEAT heatid="360" number="4" order="4" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT><EVENT eventid="34" gender="M" number="34" order="34" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="700"/><SWIMSTYLE distance="200" name="200m Schmetterling Männer" relaycount="1" stroke="FLY"/><AGEGROUPS><AGEGROUP agegroupid="340001" agemax="11" agemin="11" gender="M" name="Jahrgang 2014"><RANKINGS/></AGEGROUP><AGEGROUP agegroupid="340002" agemax="12" agemin="12" gender="M" name="Jahrgang 2013"><RANKINGS><RANKING place="1" resultid="2683"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="340003" agemax="13" agemin="13" gender="M" name="Jahrgang 2012"><RANKINGS><RANKING place="2" resultid="2684"/><RANKING place="1" resultid="2686"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="340004" agemax="14" agemin="14" gender="M" name="Jahrgang 2011"><RANKINGS><RANKING place="1" resultid="2689"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="340005" agemax="15" agemin="15" gender="M" name="Jahrgang 2010"><RANKINGS><RANKING place="1" resultid="2685"/><RANKING place="4" resultid="2687"/><RANKING place="5" resultid="2688"/><RANKING place="2" resultid="2690"/><RANKING place="3" resultid="2694"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="340006" agemax="16" agemin="16" gender="M" name="Jahrgang 2009"><RANKINGS><RANKING place="2" resultid="2691"/><RANKING place="1" resultid="2693"/><RANKING place="3" resultid="2695"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="340007" agemax="17" agemin="17" gender="M" name="Jahrgang 2008"><RANKINGS><RANKING place="1" resultid="2692"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="340008" agemax="-1" agemin="18" gender="M" name="Jahrgang 2007 und älter"><RANKINGS/></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="361" number="1" order="1" status="OFFICIAL"/><HEAT heatid="362" number="2" order="2" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT></EVENTS></SESSION><SESSION course="LCM" date="2025-03-16" daytime="14:00" name="Abschnitt 5" number="5" warmupfrom="13:00" warmupuntil="14:00"><POOL name="Erlangen" lanemax="8" lanemin="1" type="INDOOR"/><JUDGES/><EVENTS><EVENT eventid="35" gender="F" number="35" order="35" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="700"/><SWIMSTYLE distance="50" name="50m Schmetterling Frauen" relaycount="1" stroke="FLY"/><AGEGROUPS><AGEGROUP agegroupid="350001" agemax="9" agemin="9" gender="F" name="Jahrgang 2016"><RANKINGS><RANKING place="4" resultid="2703"/><RANKING place="5" resultid="2708"/><RANKING place="1" resultid="2713"/><RANKING place="2" resultid="2714"/><RANKING place="3" resultid="2725"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="350002" agemax="10" agemin="10" gender="F" name="Jahrgang 2015"><RANKINGS><RANKING place="8" resultid="2702"/><RANKING place="9" resultid="2706"/><RANKING place="10" resultid="2709"/><RANKING place="6" resultid="2710"/><RANKING place="5" resultid="2716"/><RANKING place="7" resultid="2718"/><RANKING place="1" resultid="2721"/><RANKING place="4" resultid="2734"/><RANKING place="3" resultid="2737"/><RANKING place="2" resultid="2738"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="350003" agemax="11" agemin="11" gender="F" name="Jahrgang 2014"><RANKINGS><RANKING place="-1" resultid="2698"/><RANKING place="16" resultid="2699"/><RANKING place="17" resultid="2701"/><RANKING place="18" resultid="2704"/><RANKING place="13" resultid="2705"/><RANKING place="15" resultid="2707"/><RANKING place="14" resultid="2711"/><RANKING place="7" resultid="2712"/><RANKING place="9" resultid="2715"/><RANKING place="12" resultid="2717"/><RANKING place="11" resultid="2719"/><RANKING place="10" resultid="2722"/><RANKING place="3" resultid="2723"/><RANKING place="8" resultid="2724"/><RANKING place="4" resultid="2735"/><RANKING place="6" resultid="2740"/><RANKING place="1" resultid="2745"/><RANKING place="5" resultid="2749"/><RANKING place="2" resultid="2766"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="350004" agemax="12" agemin="12" gender="F" name="Jahrgang 2013"><RANKINGS><RANKING place="13" resultid="2696"/><RANKING place="15" resultid="2697"/><RANKING place="14" resultid="2700"/><RANKING place="12" resultid="2726"/><RANKING place="10" resultid="2729"/><RANKING place="7" resultid="2730"/><RANKING place="-1" resultid="2733"/><RANKING place="9" resultid="2741"/><RANKING place="11" resultid="2742"/><RANKING place="5" resultid="2746"/><RANKING place="8" resultid="2747"/><RANKING place="-1" resultid="2753"/><RANKING place="6" resultid="2757"/><RANKING place="4" resultid="2769"/><RANKING place="3" resultid="2771"/><RANKING place="1" resultid="2778"/><RANKING place="2" resultid="2781"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="350005" agemax="13" agemin="13" gender="F" name="Jahrgang 2012"><RANKINGS><RANKING place="19" resultid="2732"/><RANKING place="13" resultid="2736"/><RANKING place="18" resultid="2744"/><RANKING place="15" resultid="2754"/><RANKING place="16" resultid="2755"/><RANKING place="17" resultid="2759"/><RANKING place="14" resultid="2767"/><RANKING place="7" resultid="2773"/><RANKING place="8" resultid="2774"/><RANKING place="10" resultid="2776"/><RANKING place="12" resultid="2780"/><RANKING place="5" resultid="2790"/><RANKING place="4" resultid="2791"/><RANKING place="11" resultid="2796"/><RANKING place="6" resultid="2797"/><RANKING place="2" resultid="2798"/><RANKING place="9" resultid="2811"/><RANKING place="3" resultid="2818"/><RANKING place="1" resultid="2825"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="350006" agemax="14" agemin="14" gender="F" name="Jahrgang 2011"><RANKINGS><RANKING place="24" resultid="2727"/><RANKING place="22" resultid="2728"/><RANKING place="23" resultid="2731"/><RANKING place="18" resultid="2751"/><RANKING place="14" resultid="2752"/><RANKING place="19" resultid="2760"/><RANKING place="16" resultid="2761"/><RANKING place="21" resultid="2764"/><RANKING place="20" resultid="2765"/><RANKING place="17" resultid="2772"/><RANKING place="-1" resultid="2785"/><RANKING place="11" resultid="2786"/><RANKING place="10" resultid="2793"/><RANKING place="7" resultid="2794"/><RANKING place="15" resultid="2799"/><RANKING place="4" resultid="2806"/><RANKING place="3" resultid="2807"/><RANKING place="9" resultid="2809"/><RANKING place="5" resultid="2815"/><RANKING place="13" resultid="2821"/><RANKING place="12" resultid="2826"/><RANKING place="6" resultid="2835"/><RANKING place="2" resultid="2837"/><RANKING place="8" resultid="2840"/><RANKING place="1" resultid="2845"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="350007" agemax="15" agemin="15" gender="F" name="Jahrgang 2010"><RANKINGS><RANKING place="11" resultid="2739"/><RANKING place="14" resultid="2748"/><RANKING place="13" resultid="2756"/><RANKING place="12" resultid="2758"/><RANKING place="10" resultid="2762"/><RANKING place="8" resultid="2770"/><RANKING place="7" resultid="2775"/><RANKING place="9" resultid="2787"/><RANKING place="6" resultid="2792"/><RANKING place="3" resultid="2812"/><RANKING place="5" resultid="2819"/><RANKING place="4" resultid="2820"/><RANKING place="2" resultid="2833"/><RANKING place="1" resultid="2851"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="350008" agemax="16" agemin="16" gender="F" name="Jahrgang 2009"><RANKINGS><RANKING place="19" resultid="2743"/><RANKING place="-1" resultid="2750"/><RANKING place="15" resultid="2763"/><RANKING place="18" resultid="2768"/><RANKING place="11" resultid="2779"/><RANKING place="17" resultid="2782"/><RANKING place="14" resultid="2784"/><RANKING place="16" resultid="2789"/><RANKING place="10" resultid="2800"/><RANKING place="8" resultid="2801"/><RANKING place="12" resultid="2803"/><RANKING place="9" resultid="2804"/><RANKING place="13" resultid="2805"/><RANKING place="-1" resultid="2808"/><RANKING place="-1" resultid="2810"/><RANKING place="7" resultid="2816"/><RANKING place="4" resultid="2823"/><RANKING place="5" resultid="2824"/><RANKING place="-1" resultid="2827"/><RANKING place="6" resultid="2828"/><RANKING place="3" resultid="2841"/><RANKING place="2" resultid="2844"/><RANKING place="1" resultid="2847"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="350009" agemax="17" agemin="17" gender="F" name="Jahrgang 2008"><RANKINGS><RANKING place="6" resultid="2788"/><RANKING place="5" resultid="2795"/><RANKING place="4" resultid="2802"/><RANKING place="2" resultid="2813"/><RANKING place="-1" resultid="2829"/><RANKING place="1" resultid="2831"/><RANKING place="3" resultid="2839"/><RANKING place="-1" resultid="2843"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="350010" agemax="-1" agemin="18" gender="F" name="Jahrgang 2007 und älter"><RANKINGS><RANKING place="15" resultid="2720"/><RANKING place="12" resultid="2777"/><RANKING place="14" resultid="2783"/><RANKING place="-1" resultid="2814"/><RANKING place="13" resultid="2817"/><RANKING place="9" resultid="2822"/><RANKING place="8" resultid="2830"/><RANKING place="6" resultid="2832"/><RANKING place="10" resultid="2834"/><RANKING place="11" resultid="2836"/><RANKING place="5" resultid="2838"/><RANKING place="7" resultid="2842"/><RANKING place="2" resultid="2846"/><RANKING place="1" resultid="2848"/><RANKING place="3" resultid="2849"/><RANKING place="4" resultid="2850"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="363" number="1" order="1" status="OFFICIAL"/><HEAT heatid="364" number="2" order="2" status="OFFICIAL"/><HEAT heatid="365" number="3" order="3" status="OFFICIAL"/><HEAT heatid="366" number="4" order="4" status="OFFICIAL"/><HEAT heatid="367" number="5" order="5" status="OFFICIAL"/><HEAT heatid="368" number="6" order="6" status="OFFICIAL"/><HEAT heatid="369" number="7" order="7" status="OFFICIAL"/><HEAT heatid="370" number="8" order="8" status="OFFICIAL"/><HEAT heatid="371" number="9" order="9" status="OFFICIAL"/><HEAT heatid="372" number="10" order="10" status="OFFICIAL"/><HEAT heatid="373" number="11" order="11" status="OFFICIAL"/><HEAT heatid="374" number="12" order="12" status="OFFICIAL"/><HEAT heatid="375" number="13" order="13" status="OFFICIAL"/><HEAT heatid="376" number="14" order="14" status="OFFICIAL"/><HEAT heatid="377" number="15" order="15" status="OFFICIAL"/><HEAT heatid="378" number="16" order="16" status="OFFICIAL"/><HEAT heatid="379" number="17" order="17" status="OFFICIAL"/><HEAT heatid="380" number="18" order="18" status="OFFICIAL"/><HEAT heatid="381" number="19" order="19" status="OFFICIAL"/><HEAT heatid="382" number="20" order="20" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT><EVENT eventid="36" gender="M" number="36" order="36" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="700"/><SWIMSTYLE distance="50" name="50m Schmetterling Männer" relaycount="1" stroke="FLY"/><AGEGROUPS><AGEGROUP agegroupid="360001" agemax="9" agemin="9" gender="M" name="Jahrgang 2016"><RANKINGS><RANKING place="1" resultid="2852"/><RANKING place="2" resultid="2861"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="360002" agemax="10" agemin="10" gender="M" name="Jahrgang 2015"><RANKINGS><RANKING place="12" resultid="2854"/><RANKING place="6" resultid="2857"/><RANKING place="11" resultid="2860"/><RANKING place="10" resultid="2863"/><RANKING place="9" resultid="2869"/><RANKING place="5" resultid="2874"/><RANKING place="8" resultid="2876"/><RANKING place="7" resultid="2884"/><RANKING place="1" resultid="2886"/><RANKING place="3" resultid="2887"/><RANKING place="3" resultid="2890"/><RANKING place="2" resultid="2892"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="360003" agemax="11" agemin="11" gender="M" name="Jahrgang 2014"><RANKINGS><RANKING place="-1" resultid="2856"/><RANKING place="7" resultid="2858"/><RANKING place="9" resultid="2865"/><RANKING place="6" resultid="2870"/><RANKING place="8" resultid="2880"/><RANKING place="5" resultid="2885"/><RANKING place="2" resultid="2888"/><RANKING place="1" resultid="2893"/><RANKING place="4" resultid="2900"/><RANKING place="3" resultid="2901"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="360004" agemax="12" agemin="12" gender="M" name="Jahrgang 2013"><RANKINGS><RANKING place="11" resultid="2853"/><RANKING place="-1" resultid="2855"/><RANKING place="13" resultid="2859"/><RANKING place="-1" resultid="2862"/><RANKING place="5" resultid="2864"/><RANKING place="4" resultid="2866"/><RANKING place="3" resultid="2867"/><RANKING place="8" resultid="2872"/><RANKING place="9" resultid="2873"/><RANKING place="10" resultid="2875"/><RANKING place="12" resultid="2877"/><RANKING place="6" resultid="2878"/><RANKING place="7" resultid="2881"/><RANKING place="2" resultid="2894"/><RANKING place="1" resultid="2917"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="360005" agemax="13" agemin="13" gender="M" name="Jahrgang 2012"><RANKINGS><RANKING place="10" resultid="2868"/><RANKING place="-1" resultid="2871"/><RANKING place="11" resultid="2879"/><RANKING place="8" resultid="2889"/><RANKING place="5" resultid="2899"/><RANKING place="6" resultid="2906"/><RANKING place="3" resultid="2907"/><RANKING place="9" resultid="2908"/><RANKING place="7" resultid="2911"/><RANKING place="4" resultid="2914"/><RANKING place="1" resultid="2923"/><RANKING place="2" resultid="2941"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="360006" agemax="14" agemin="14" gender="M" name="Jahrgang 2011"><RANKINGS><RANKING place="-1" resultid="2883"/><RANKING place="15" resultid="2891"/><RANKING place="10" resultid="2895"/><RANKING place="18" resultid="2896"/><RANKING place="19" resultid="2898"/><RANKING place="17" resultid="2902"/><RANKING place="12" resultid="2905"/><RANKING place="14" resultid="2909"/><RANKING place="11" resultid="2910"/><RANKING place="9" resultid="2913"/><RANKING place="-1" resultid="2920"/><RANKING place="8" resultid="2921"/><RANKING place="16" resultid="2924"/><RANKING place="1" resultid="2931"/><RANKING place="7" resultid="2932"/><RANKING place="13" resultid="2933"/><RANKING place="4" resultid="2936"/><RANKING place="6" resultid="2939"/><RANKING place="5" resultid="2942"/><RANKING place="2" resultid="2956"/><RANKING place="3" resultid="2957"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="360007" agemax="15" agemin="15" gender="M" name="Jahrgang 2010"><RANKINGS><RANKING place="17" resultid="2897"/><RANKING place="15" resultid="2904"/><RANKING place="13" resultid="2912"/><RANKING place="20" resultid="2915"/><RANKING place="14" resultid="2916"/><RANKING place="16" resultid="2918"/><RANKING place="18" resultid="2922"/><RANKING place="19" resultid="2925"/><RANKING place="11" resultid="2926"/><RANKING place="9" resultid="2929"/><RANKING place="10" resultid="2930"/><RANKING place="12" resultid="2940"/><RANKING place="7" resultid="2943"/><RANKING place="8" resultid="2949"/><RANKING place="6" resultid="2950"/><RANKING place="5" resultid="2959"/><RANKING place="4" resultid="2961"/><RANKING place="2" resultid="2969"/><RANKING place="3" resultid="2970"/><RANKING place="1" resultid="2983"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="360008" agemax="16" agemin="16" gender="M" name="Jahrgang 2009"><RANKINGS><RANKING place="19" resultid="2919"/><RANKING place="16" resultid="2927"/><RANKING place="18" resultid="2935"/><RANKING place="12" resultid="2937"/><RANKING place="17" resultid="2938"/><RANKING place="-1" resultid="2946"/><RANKING place="15" resultid="2947"/><RANKING place="8" resultid="2948"/><RANKING place="14" resultid="2951"/><RANKING place="10" resultid="2952"/><RANKING place="13" resultid="2953"/><RANKING place="9" resultid="2958"/><RANKING place="11" resultid="2965"/><RANKING place="3" resultid="2972"/><RANKING place="7" resultid="2973"/><RANKING place="4" resultid="2974"/><RANKING place="6" resultid="2975"/><RANKING place="5" resultid="2976"/><RANKING place="1" resultid="2979"/><RANKING place="2" resultid="2988"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="360009" agemax="17" agemin="17" gender="M" name="Jahrgang 2008"><RANKINGS><RANKING place="7" resultid="2882"/><RANKING place="8" resultid="2928"/><RANKING place="9" resultid="2934"/><RANKING place="6" resultid="2945"/><RANKING place="-1" resultid="2960"/><RANKING place="4" resultid="2962"/><RANKING place="5" resultid="2964"/><RANKING place="-1" resultid="2981"/><RANKING place="1" resultid="2984"/><RANKING place="2" resultid="2985"/><RANKING place="3" resultid="2987"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="360010" agemax="-1" agemin="18" gender="M" name="Jahrgang 2007 und älter"><RANKINGS><RANKING place="13" resultid="2903"/><RANKING place="11" resultid="2944"/><RANKING place="7" resultid="2954"/><RANKING place="12" resultid="2955"/><RANKING place="9" resultid="2963"/><RANKING place="10" resultid="2966"/><RANKING place="6" resultid="2967"/><RANKING place="-1" resultid="2968"/><RANKING place="8" resultid="2971"/><RANKING place="2" resultid="2977"/><RANKING place="4" resultid="2978"/><RANKING place="3" resultid="2980"/><RANKING place="1" resultid="2982"/><RANKING place="5" resultid="2986"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="383" number="1" order="1" status="OFFICIAL"/><HEAT heatid="384" number="2" order="2" status="OFFICIAL"/><HEAT heatid="385" number="3" order="3" status="OFFICIAL"/><HEAT heatid="386" number="4" order="4" status="OFFICIAL"/><HEAT heatid="387" number="5" order="5" status="OFFICIAL"/><HEAT heatid="388" number="6" order="6" status="OFFICIAL"/><HEAT heatid="389" number="7" order="7" status="OFFICIAL"/><HEAT heatid="390" number="8" order="8" status="OFFICIAL"/><HEAT heatid="391" number="9" order="9" status="OFFICIAL"/><HEAT heatid="392" number="10" order="10" status="OFFICIAL"/><HEAT heatid="393" number="11" order="11" status="OFFICIAL"/><HEAT heatid="394" number="12" order="12" status="OFFICIAL"/><HEAT heatid="395" number="13" order="13" status="OFFICIAL"/><HEAT heatid="396" number="14" order="14" status="OFFICIAL"/><HEAT heatid="397" number="15" order="15" status="OFFICIAL"/><HEAT heatid="398" number="16" order="16" status="OFFICIAL"/><HEAT heatid="399" number="17" order="17" status="OFFICIAL"/><HEAT heatid="400" number="18" order="18" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT><EVENT eventid="37" gender="F" number="37" order="37" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="700"/><SWIMSTYLE distance="200" name="200m Rücken Frauen" relaycount="1" stroke="BACK"/><AGEGROUPS><AGEGROUP agegroupid="370001" agemax="9" agemin="9" gender="F" name="Jahrgang 2016"><RANKINGS><RANKING place="-1" resultid="2990"/><RANKING place="4" resultid="2997"/><RANKING place="3" resultid="3001"/><RANKING place="2" resultid="3004"/><RANKING place="1" resultid="3005"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="370002" agemax="10" agemin="10" gender="F" name="Jahrgang 2015"><RANKINGS><RANKING place="7" resultid="2989"/><RANKING place="6" resultid="2991"/><RANKING place="5" resultid="2992"/><RANKING place="4" resultid="2996"/><RANKING place="3" resultid="2998"/><RANKING place="1" resultid="3007"/><RANKING place="2" resultid="3015"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="370003" agemax="11" agemin="11" gender="F" name="Jahrgang 2014"><RANKINGS><RANKING place="8" resultid="2993"/><RANKING place="9" resultid="2994"/><RANKING place="-1" resultid="2999"/><RANKING place="-1" resultid="3000"/><RANKING place="7" resultid="3002"/><RANKING place="11" resultid="3003"/><RANKING place="6" resultid="3006"/><RANKING place="10" resultid="3010"/><RANKING place="5" resultid="3012"/><RANKING place="4" resultid="3020"/><RANKING place="2" resultid="3025"/><RANKING place="1" resultid="3026"/><RANKING place="3" resultid="3034"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="370004" agemax="12" agemin="12" gender="F" name="Jahrgang 2013"><RANKINGS><RANKING place="13" resultid="2995"/><RANKING place="14" resultid="3009"/><RANKING place="11" resultid="3011"/><RANKING place="12" resultid="3013"/><RANKING place="-1" resultid="3019"/><RANKING place="10" resultid="3021"/><RANKING place="9" resultid="3022"/><RANKING place="6" resultid="3024"/><RANKING place="5" resultid="3028"/><RANKING place="8" resultid="3029"/><RANKING place="7" resultid="3030"/><RANKING place="3" resultid="3033"/><RANKING place="4" resultid="3036"/><RANKING place="-1" resultid="3039"/><RANKING place="2" resultid="3047"/><RANKING place="1" resultid="3060"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="370005" agemax="13" agemin="13" gender="F" name="Jahrgang 2012"><RANKINGS><RANKING place="8" resultid="3014"/><RANKING place="7" resultid="3016"/><RANKING place="6" resultid="3017"/><RANKING place="4" resultid="3023"/><RANKING place="5" resultid="3027"/><RANKING place="3" resultid="3044"/><RANKING place="2" resultid="3069"/><RANKING place="1" resultid="3070"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="370006" agemax="14" agemin="14" gender="F" name="Jahrgang 2011"><RANKINGS><RANKING place="10" resultid="3035"/><RANKING place="8" resultid="3040"/><RANKING place="9" resultid="3041"/><RANKING place="5" resultid="3048"/><RANKING place="3" resultid="3053"/><RANKING place="11" resultid="3054"/><RANKING place="7" resultid="3055"/><RANKING place="6" resultid="3058"/><RANKING place="4" resultid="3059"/><RANKING place="2" resultid="3065"/><RANKING place="1" resultid="3072"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="370007" agemax="15" agemin="15" gender="F" name="Jahrgang 2010"><RANKINGS><RANKING place="9" resultid="3018"/><RANKING place="-1" resultid="3032"/><RANKING place="8" resultid="3038"/><RANKING place="7" resultid="3045"/><RANKING place="4" resultid="3049"/><RANKING place="5" resultid="3050"/><RANKING place="3" resultid="3063"/><RANKING place="6" resultid="3064"/><RANKING place="2" resultid="3071"/><RANKING place="1" resultid="3077"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="370008" agemax="16" agemin="16" gender="F" name="Jahrgang 2009"><RANKINGS><RANKING place="11" resultid="3008"/><RANKING place="9" resultid="3031"/><RANKING place="10" resultid="3046"/><RANKING place="7" resultid="3051"/><RANKING place="8" resultid="3052"/><RANKING place="6" resultid="3056"/><RANKING place="5" resultid="3061"/><RANKING place="-1" resultid="3067"/><RANKING place="2" resultid="3068"/><RANKING place="4" resultid="3074"/><RANKING place="1" resultid="3075"/><RANKING place="3" resultid="3076"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="370009" agemax="17" agemin="17" gender="F" name="Jahrgang 2008"><RANKINGS><RANKING place="1" resultid="3057"/><RANKING place="2" resultid="3062"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="370010" agemax="-1" agemin="18" gender="F" name="Jahrgang 2007 und älter"><RANKINGS><RANKING place="5" resultid="3037"/><RANKING place="3" resultid="3042"/><RANKING place="4" resultid="3043"/><RANKING place="2" resultid="3066"/><RANKING place="1" resultid="3073"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="401" number="1" order="1" status="OFFICIAL"/><HEAT heatid="402" number="2" order="2" status="OFFICIAL"/><HEAT heatid="403" number="3" order="3" status="OFFICIAL"/><HEAT heatid="404" number="4" order="4" status="OFFICIAL"/><HEAT heatid="405" number="5" order="5" status="OFFICIAL"/><HEAT heatid="406" number="6" order="6" status="OFFICIAL"/><HEAT heatid="407" number="7" order="7" status="OFFICIAL"/><HEAT heatid="408" number="8" order="8" status="OFFICIAL"/><HEAT heatid="409" number="9" order="9" status="OFFICIAL"/><HEAT heatid="410" number="10" order="10" status="OFFICIAL"/><HEAT heatid="411" number="11" order="11" status="OFFICIAL"/><HEAT heatid="412" number="12" order="12" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT><EVENT eventid="38" gender="M" number="38" order="38" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="700"/><SWIMSTYLE distance="200" name="200m Rücken Männer" relaycount="1" stroke="BACK"/><AGEGROUPS><AGEGROUP agegroupid="380001" agemax="9" agemin="9" gender="M" name="Jahrgang 2016"><RANKINGS><RANKING place="2" resultid="3079"/><RANKING place="1" resultid="3088"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="380002" agemax="10" agemin="10" gender="M" name="Jahrgang 2015"><RANKINGS><RANKING place="-1" resultid="3080"/><RANKING place="-1" resultid="3081"/><RANKING place="8" resultid="3083"/><RANKING place="1" resultid="3087"/><RANKING place="7" resultid="3089"/><RANKING place="-1" resultid="3090"/><RANKING place="3" resultid="3091"/><RANKING place="6" resultid="3092"/><RANKING place="4" resultid="3096"/><RANKING place="2" resultid="3097"/><RANKING place="5" resultid="3098"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="380003" agemax="11" agemin="11" gender="M" name="Jahrgang 2014"><RANKINGS><RANKING place="6" resultid="3078"/><RANKING place="7" resultid="3084"/><RANKING place="4" resultid="3085"/><RANKING place="2" resultid="3093"/><RANKING place="3" resultid="3094"/><RANKING place="5" resultid="3095"/><RANKING place="1" resultid="3103"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="380004" agemax="12" agemin="12" gender="M" name="Jahrgang 2013"><RANKINGS><RANKING place="5" resultid="3082"/><RANKING place="7" resultid="3086"/><RANKING place="3" resultid="3099"/><RANKING place="6" resultid="3101"/><RANKING place="4" resultid="3102"/><RANKING place="1" resultid="3109"/><RANKING place="2" resultid="3120"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="380005" agemax="13" agemin="13" gender="M" name="Jahrgang 2012"><RANKINGS><RANKING place="1" resultid="3111"/><RANKING place="3" resultid="3112"/><RANKING place="2" resultid="3114"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="380006" agemax="14" agemin="14" gender="M" name="Jahrgang 2011"><RANKINGS><RANKING place="4" resultid="3100"/><RANKING place="6" resultid="3105"/><RANKING place="5" resultid="3106"/><RANKING place="2" resultid="3108"/><RANKING place="3" resultid="3110"/><RANKING place="-1" resultid="3113"/><RANKING place="-1" resultid="3115"/><RANKING place="1" resultid="3118"/><RANKING place="-1" resultid="3119"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="380007" agemax="15" agemin="15" gender="M" name="Jahrgang 2010"><RANKINGS><RANKING place="4" resultid="3104"/><RANKING place="3" resultid="3116"/><RANKING place="2" resultid="3121"/><RANKING place="1" resultid="3125"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="380008" agemax="16" agemin="16" gender="M" name="Jahrgang 2009"><RANKINGS><RANKING place="3" resultid="3107"/><RANKING place="1" resultid="3123"/><RANKING place="2" resultid="3126"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="380009" agemax="17" agemin="17" gender="M" name="Jahrgang 2008"><RANKINGS><RANKING place="1" resultid="3122"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="380010" agemax="-1" agemin="18" gender="M" name="Jahrgang 2007 und älter"><RANKINGS><RANKING place="-1" resultid="3117"/><RANKING place="1" resultid="3124"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="413" number="1" order="1" status="OFFICIAL"/><HEAT heatid="414" number="2" order="2" status="OFFICIAL"/><HEAT heatid="415" number="3" order="3" status="OFFICIAL"/><HEAT heatid="416" number="4" order="4" status="OFFICIAL"/><HEAT heatid="417" number="5" order="5" status="OFFICIAL"/><HEAT heatid="418" number="6" order="6" status="OFFICIAL"/><HEAT heatid="419" number="7" order="7" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT><EVENT eventid="39" gender="F" number="39" order="39" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="700"/><SWIMSTYLE distance="100" name="100m Freistil Frauen" relaycount="1" stroke="FREE"/><AGEGROUPS><AGEGROUP agegroupid="390001" agemax="8" agemin="8" gender="F" name="Jahrgang 2017"><RANKINGS><RANKING place="2" resultid="3131"/><RANKING place="4" resultid="3137"/><RANKING place="3" resultid="3140"/><RANKING place="5" resultid="3141"/><RANKING place="1" resultid="3160"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="390002" agemax="9" agemin="9" gender="F" name="Jahrgang 2016"><RANKINGS><RANKING place="12" resultid="3128"/><RANKING place="13" resultid="3138"/><RANKING place="11" resultid="3139"/><RANKING place="10" resultid="3145"/><RANKING place="6" resultid="3157"/><RANKING place="9" resultid="3165"/><RANKING place="8" resultid="3170"/><RANKING place="5" resultid="3172"/><RANKING place="7" resultid="3176"/><RANKING place="4" resultid="3179"/><RANKING place="3" resultid="3200"/><RANKING place="2" resultid="3202"/><RANKING place="1" resultid="3203"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="390003" agemax="10" agemin="10" gender="F" name="Jahrgang 2015"><RANKINGS><RANKING place="24" resultid="3129"/><RANKING place="18" resultid="3135"/><RANKING place="21" resultid="3136"/><RANKING place="23" resultid="3143"/><RANKING place="22" resultid="3144"/><RANKING place="20" resultid="3146"/><RANKING place="13" resultid="3149"/><RANKING place="14" resultid="3151"/><RANKING place="16" resultid="3153"/><RANKING place="19" resultid="3161"/><RANKING place="12" resultid="3167"/><RANKING place="17" resultid="3171"/><RANKING place="4" resultid="3174"/><RANKING place="3" resultid="3175"/><RANKING place="9" resultid="3180"/><RANKING place="-1" resultid="3182"/><RANKING place="10" resultid="3183"/><RANKING place="8" resultid="3184"/><RANKING place="15" resultid="3185"/><RANKING place="6" resultid="3187"/><RANKING place="11" resultid="3192"/><RANKING place="5" resultid="3194"/><RANKING place="7" resultid="3201"/><RANKING place="2" resultid="3233"/><RANKING place="1" resultid="3234"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="390004" agemax="11" agemin="11" gender="F" name="Jahrgang 2014"><RANKINGS><RANKING place="29" resultid="3127"/><RANKING place="32" resultid="3132"/><RANKING place="34" resultid="3134"/><RANKING place="27" resultid="3147"/><RANKING place="35" resultid="3148"/><RANKING place="31" resultid="3150"/><RANKING place="30" resultid="3152"/><RANKING place="28" resultid="3154"/><RANKING place="26" resultid="3156"/><RANKING place="33" resultid="3162"/><RANKING place="24" resultid="3168"/><RANKING place="23" resultid="3169"/><RANKING place="-1" resultid="3177"/><RANKING place="22" resultid="3181"/><RANKING place="11" resultid="3186"/><RANKING place="20" resultid="3188"/><RANKING place="18" resultid="3189"/><RANKING place="21" resultid="3190"/><RANKING place="12" resultid="3191"/><RANKING place="13" resultid="3193"/><RANKING place="15" resultid="3199"/><RANKING place="19" resultid="3204"/><RANKING place="25" resultid="3209"/><RANKING place="14" resultid="3210"/><RANKING place="9" resultid="3215"/><RANKING place="16" resultid="3216"/><RANKING place="17" resultid="3217"/><RANKING place="7" resultid="3219"/><RANKING place="10" resultid="3220"/><RANKING place="-1" resultid="3221"/><RANKING place="5" resultid="3236"/><RANKING place="8" resultid="3237"/><RANKING place="4" resultid="3239"/><RANKING place="1" resultid="3244"/><RANKING place="6" resultid="3249"/><RANKING place="3" resultid="3255"/><RANKING place="2" resultid="3267"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="390005" agemax="12" agemin="12" gender="F" name="Jahrgang 2013"><RANKINGS><RANKING place="30" resultid="3130"/><RANKING place="25" resultid="3133"/><RANKING place="28" resultid="3142"/><RANKING place="24" resultid="3155"/><RANKING place="27" resultid="3158"/><RANKING place="23" resultid="3159"/><RANKING place="19" resultid="3163"/><RANKING place="29" resultid="3164"/><RANKING place="26" resultid="3166"/><RANKING place="-1" resultid="3173"/><RANKING place="20" resultid="3195"/><RANKING place="21" resultid="3196"/><RANKING place="22" resultid="3198"/><RANKING place="18" resultid="3208"/><RANKING place="15" resultid="3211"/><RANKING place="16" resultid="3212"/><RANKING place="-1" resultid="3224"/><RANKING place="8" resultid="3228"/><RANKING place="7" resultid="3230"/><RANKING place="12" resultid="3231"/><RANKING place="17" resultid="3232"/><RANKING place="11" resultid="3242"/><RANKING place="13" resultid="3245"/><RANKING place="10" resultid="3252"/><RANKING place="9" resultid="3256"/><RANKING place="14" resultid="3257"/><RANKING place="6" resultid="3258"/><RANKING place="-1" resultid="3259"/><RANKING place="5" resultid="3261"/><RANKING place="4" resultid="3272"/><RANKING place="2" resultid="3282"/><RANKING place="3" resultid="3284"/><RANKING place="1" resultid="3318"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="390006" agemax="13" agemin="13" gender="F" name="Jahrgang 2012"><RANKINGS><RANKING place="18" resultid="3197"/><RANKING place="17" resultid="3205"/><RANKING place="15" resultid="3214"/><RANKING place="-1" resultid="3222"/><RANKING place="13" resultid="3235"/><RANKING place="16" resultid="3246"/><RANKING place="10" resultid="3253"/><RANKING place="14" resultid="3254"/><RANKING place="12" resultid="3263"/><RANKING place="8" resultid="3277"/><RANKING place="11" resultid="3280"/><RANKING place="3" resultid="3283"/><RANKING place="5" resultid="3292"/><RANKING place="7" resultid="3294"/><RANKING place="9" resultid="3301"/><RANKING place="6" resultid="3312"/><RANKING place="2" resultid="3325"/><RANKING place="4" resultid="3328"/><RANKING place="1" resultid="3348"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="390007" agemax="14" agemin="14" gender="F" name="Jahrgang 2011"><RANKINGS><RANKING place="28" resultid="3206"/><RANKING place="26" resultid="3213"/><RANKING place="27" resultid="3218"/><RANKING place="23" resultid="3225"/><RANKING place="19" resultid="3238"/><RANKING place="24" resultid="3240"/><RANKING place="25" resultid="3250"/><RANKING place="-1" resultid="3262"/><RANKING place="20" resultid="3266"/><RANKING place="14" resultid="3268"/><RANKING place="11" resultid="3279"/><RANKING place="-1" resultid="3288"/><RANKING place="21" resultid="3290"/><RANKING place="18" resultid="3295"/><RANKING place="3" resultid="3298"/><RANKING place="17" resultid="3302"/><RANKING place="13" resultid="3304"/><RANKING place="6" resultid="3306"/><RANKING place="8" resultid="3307"/><RANKING place="22" resultid="3311"/><RANKING place="15" resultid="3315"/><RANKING place="16" resultid="3319"/><RANKING place="10" resultid="3322"/><RANKING place="5" resultid="3323"/><RANKING place="1" resultid="3324"/><RANKING place="12" resultid="3331"/><RANKING place="4" resultid="3332"/><RANKING place="7" resultid="3337"/><RANKING place="9" resultid="3340"/><RANKING place="2" resultid="3344"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="390008" agemax="15" agemin="15" gender="F" name="Jahrgang 2010"><RANKINGS><RANKING place="22" resultid="3223"/><RANKING place="21" resultid="3226"/><RANKING place="19" resultid="3248"/><RANKING place="16" resultid="3265"/><RANKING place="20" resultid="3270"/><RANKING place="-1" resultid="3271"/><RANKING place="18" resultid="3273"/><RANKING place="17" resultid="3276"/><RANKING place="15" resultid="3281"/><RANKING place="14" resultid="3287"/><RANKING place="9" resultid="3291"/><RANKING place="11" resultid="3293"/><RANKING place="13" resultid="3296"/><RANKING place="10" resultid="3299"/><RANKING place="8" resultid="3303"/><RANKING place="12" resultid="3320"/><RANKING place="7" resultid="3326"/><RANKING place="5" resultid="3342"/><RANKING place="6" resultid="3345"/><RANKING place="4" resultid="3347"/><RANKING place="3" resultid="3352"/><RANKING place="2" resultid="3354"/><RANKING place="1" resultid="3362"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="390009" agemax="16" agemin="16" gender="F" name="Jahrgang 2009"><RANKINGS><RANKING place="25" resultid="3178"/><RANKING place="-1" resultid="3227"/><RANKING place="19" resultid="3229"/><RANKING place="24" resultid="3241"/><RANKING place="21" resultid="3243"/><RANKING place="22" resultid="3251"/><RANKING place="20" resultid="3260"/><RANKING place="23" resultid="3264"/><RANKING place="17" resultid="3275"/><RANKING place="18" resultid="3278"/><RANKING place="8" resultid="3285"/><RANKING place="16" resultid="3297"/><RANKING place="13" resultid="3308"/><RANKING place="10" resultid="3313"/><RANKING place="14" resultid="3314"/><RANKING place="12" resultid="3316"/><RANKING place="15" resultid="3317"/><RANKING place="11" resultid="3321"/><RANKING place="-1" resultid="3327"/><RANKING place="9" resultid="3329"/><RANKING place="7" resultid="3333"/><RANKING place="6" resultid="3335"/><RANKING place="5" resultid="3338"/><RANKING place="4" resultid="3346"/><RANKING place="-1" resultid="3351"/><RANKING place="1" resultid="3355"/><RANKING place="2" resultid="3356"/><RANKING place="3" resultid="3357"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="390010" agemax="17" agemin="17" gender="F" name="Jahrgang 2008"><RANKINGS><RANKING place="5" resultid="3289"/><RANKING place="3" resultid="3336"/><RANKING place="4" resultid="3341"/><RANKING place="-1" resultid="3350"/><RANKING place="1" resultid="3358"/><RANKING place="2" resultid="3360"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="390011" agemax="-1" agemin="18" gender="F" name="Jahrgang 2007 und älter"><RANKINGS><RANKING place="19" resultid="3207"/><RANKING place="18" resultid="3247"/><RANKING place="15" resultid="3269"/><RANKING place="14" resultid="3274"/><RANKING place="13" resultid="3286"/><RANKING place="17" resultid="3300"/><RANKING place="16" resultid="3305"/><RANKING place="11" resultid="3309"/><RANKING place="10" resultid="3310"/><RANKING place="12" resultid="3330"/><RANKING place="9" resultid="3334"/><RANKING place="8" resultid="3339"/><RANKING place="-1" resultid="3343"/><RANKING place="6" resultid="3349"/><RANKING place="5" resultid="3353"/><RANKING place="4" resultid="3359"/><RANKING place="1" resultid="3361"/><RANKING place="2" resultid="3363"/><RANKING place="3" resultid="3364"/><RANKING place="7" resultid="3365"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="420" number="1" order="1" status="OFFICIAL"/><HEAT heatid="421" number="2" order="2" status="OFFICIAL"/><HEAT heatid="422" number="3" order="3" status="OFFICIAL"/><HEAT heatid="423" number="4" order="4" status="OFFICIAL"/><HEAT heatid="424" number="5" order="5" status="OFFICIAL"/><HEAT heatid="425" number="6" order="6" status="OFFICIAL"/><HEAT heatid="426" number="7" order="7" status="OFFICIAL"/><HEAT heatid="427" number="8" order="8" status="OFFICIAL"/><HEAT heatid="428" number="9" order="9" status="OFFICIAL"/><HEAT heatid="429" number="10" order="10" status="OFFICIAL"/><HEAT heatid="430" number="11" order="11" status="OFFICIAL"/><HEAT heatid="431" number="12" order="12" status="OFFICIAL"/><HEAT heatid="432" number="13" order="13" status="OFFICIAL"/><HEAT heatid="433" number="14" order="14" status="OFFICIAL"/><HEAT heatid="434" number="15" order="15" status="OFFICIAL"/><HEAT heatid="435" number="16" order="16" status="OFFICIAL"/><HEAT heatid="436" number="17" order="17" status="OFFICIAL"/><HEAT heatid="437" number="18" order="18" status="OFFICIAL"/><HEAT heatid="438" number="19" order="19" status="OFFICIAL"/><HEAT heatid="439" number="20" order="20" status="OFFICIAL"/><HEAT heatid="440" number="21" order="21" status="OFFICIAL"/><HEAT heatid="441" number="22" order="22" status="OFFICIAL"/><HEAT heatid="442" number="23" order="23" status="OFFICIAL"/><HEAT heatid="443" number="24" order="24" status="OFFICIAL"/><HEAT heatid="444" number="25" order="25" status="OFFICIAL"/><HEAT heatid="445" number="26" order="26" status="OFFICIAL"/><HEAT heatid="446" number="27" order="27" status="OFFICIAL"/><HEAT heatid="447" number="28" order="28" status="OFFICIAL"/><HEAT heatid="448" number="29" order="29" status="OFFICIAL"/><HEAT heatid="449" number="30" order="30" status="OFFICIAL"/><HEAT heatid="450" number="31" order="31" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT><EVENT eventid="40" gender="M" number="40" order="40" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="700"/><SWIMSTYLE distance="100" name="100m Freistil Männer" relaycount="1" stroke="FREE"/><AGEGROUPS><AGEGROUP agegroupid="400001" agemax="8" agemin="8" gender="M" name="Jahrgang 2017"><RANKINGS><RANKING place="1" resultid="3389"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="400002" agemax="9" agemin="9" gender="M" name="Jahrgang 2016"><RANKINGS><RANKING place="6" resultid="3374"/><RANKING place="4" resultid="3376"/><RANKING place="3" resultid="3377"/><RANKING place="5" resultid="3379"/><RANKING place="1" resultid="3385"/><RANKING place="2" resultid="3395"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="400003" agemax="10" agemin="10" gender="M" name="Jahrgang 2015"><RANKINGS><RANKING place="-1" resultid="3367"/><RANKING place="19" resultid="3375"/><RANKING place="15" resultid="3378"/><RANKING place="16" resultid="3380"/><RANKING place="10" resultid="3382"/><RANKING place="-1" resultid="3383"/><RANKING place="14" resultid="3384"/><RANKING place="18" resultid="3388"/><RANKING place="13" resultid="3392"/><RANKING place="12" resultid="3393"/><RANKING place="17" resultid="3397"/><RANKING place="9" resultid="3398"/><RANKING place="4" resultid="3400"/><RANKING place="8" resultid="3407"/><RANKING place="-1" resultid="3411"/><RANKING place="6" resultid="3414"/><RANKING place="2" resultid="3417"/><RANKING place="3" resultid="3418"/><RANKING place="11" resultid="3421"/><RANKING place="7" resultid="3430"/><RANKING place="5" resultid="3440"/><RANKING place="1" resultid="3446"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="400004" agemax="11" agemin="11" gender="M" name="Jahrgang 2014"><RANKINGS><RANKING place="24" resultid="3386"/><RANKING place="26" resultid="3387"/><RANKING place="18" resultid="3390"/><RANKING place="25" resultid="3394"/><RANKING place="10" resultid="3401"/><RANKING place="19" resultid="3402"/><RANKING place="23" resultid="3403"/><RANKING place="20" resultid="3405"/><RANKING place="21" resultid="3406"/><RANKING place="22" resultid="3412"/><RANKING place="16" resultid="3413"/><RANKING place="15" resultid="3415"/><RANKING place="6" resultid="3416"/><RANKING place="17" resultid="3420"/><RANKING place="9" resultid="3426"/><RANKING place="14" resultid="3427"/><RANKING place="11" resultid="3428"/><RANKING place="13" resultid="3429"/><RANKING place="8" resultid="3433"/><RANKING place="12" resultid="3436"/><RANKING place="7" resultid="3437"/><RANKING place="4" resultid="3444"/><RANKING place="5" resultid="3452"/><RANKING place="1" resultid="3457"/><RANKING place="3" resultid="3458"/><RANKING place="2" resultid="3459"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="400005" agemax="12" agemin="12" gender="M" name="Jahrgang 2013"><RANKINGS><RANKING place="18" resultid="3368"/><RANKING place="20" resultid="3369"/><RANKING place="16" resultid="3391"/><RANKING place="-1" resultid="3396"/><RANKING place="17" resultid="3399"/><RANKING place="19" resultid="3404"/><RANKING place="14" resultid="3422"/><RANKING place="15" resultid="3423"/><RANKING place="-1" resultid="3425"/><RANKING place="10" resultid="3434"/><RANKING place="12" resultid="3438"/><RANKING place="8" resultid="3441"/><RANKING place="11" resultid="3443"/><RANKING place="9" resultid="3447"/><RANKING place="13" resultid="3448"/><RANKING place="3" resultid="3454"/><RANKING place="6" resultid="3456"/><RANKING place="5" resultid="3461"/><RANKING place="7" resultid="3466"/><RANKING place="4" resultid="3471"/><RANKING place="2" resultid="3479"/><RANKING place="1" resultid="3496"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="400006" agemax="13" agemin="13" gender="M" name="Jahrgang 2012"><RANKINGS><RANKING place="17" resultid="3366"/><RANKING place="18" resultid="3370"/><RANKING place="19" resultid="3371"/><RANKING place="16" resultid="3372"/><RANKING place="-1" resultid="3409"/><RANKING place="15" resultid="3410"/><RANKING place="14" resultid="3424"/><RANKING place="11" resultid="3435"/><RANKING place="9" resultid="3439"/><RANKING place="12" resultid="3451"/><RANKING place="7" resultid="3460"/><RANKING place="10" resultid="3464"/><RANKING place="13" resultid="3465"/><RANKING place="8" resultid="3472"/><RANKING place="6" resultid="3476"/><RANKING place="4" resultid="3477"/><RANKING place="3" resultid="3480"/><RANKING place="2" resultid="3481"/><RANKING place="5" resultid="3486"/><RANKING place="1" resultid="3506"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="400007" agemax="14" agemin="14" gender="M" name="Jahrgang 2011"><RANKINGS><RANKING place="32" resultid="3381"/><RANKING place="31" resultid="3408"/><RANKING place="30" resultid="3419"/><RANKING place="29" resultid="3431"/><RANKING place="17" resultid="3445"/><RANKING place="26" resultid="3449"/><RANKING place="-1" resultid="3450"/><RANKING place="28" resultid="3453"/><RANKING place="25" resultid="3455"/><RANKING place="12" resultid="3462"/><RANKING place="27" resultid="3463"/><RANKING place="22" resultid="3467"/><RANKING place="24" resultid="3469"/><RANKING place="21" resultid="3473"/><RANKING place="23" resultid="3474"/><RANKING place="19" resultid="3475"/><RANKING place="16" resultid="3478"/><RANKING place="20" resultid="3482"/><RANKING place="18" resultid="3485"/><RANKING place="10" resultid="3488"/><RANKING place="14" resultid="3489"/><RANKING place="15" resultid="3490"/><RANKING place="11" resultid="3493"/><RANKING place="13" resultid="3494"/><RANKING place="7" resultid="3499"/><RANKING place="8" resultid="3501"/><RANKING place="9" resultid="3504"/><RANKING place="4" resultid="3510"/><RANKING place="5" resultid="3512"/><RANKING place="6" resultid="3514"/><RANKING place="3" resultid="3530"/><RANKING place="2" resultid="3537"/><RANKING place="1" resultid="3543"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="400008" agemax="15" agemin="15" gender="M" name="Jahrgang 2010"><RANKINGS><RANKING place="20" resultid="3373"/><RANKING place="18" resultid="3432"/><RANKING place="21" resultid="3468"/><RANKING place="16" resultid="3470"/><RANKING place="15" resultid="3483"/><RANKING place="19" resultid="3484"/><RANKING place="14" resultid="3487"/><RANKING place="17" resultid="3491"/><RANKING place="12" resultid="3492"/><RANKING place="13" resultid="3497"/><RANKING place="11" resultid="3502"/><RANKING place="10" resultid="3508"/><RANKING place="-1" resultid="3509"/><RANKING place="7" resultid="3515"/><RANKING place="8" resultid="3518"/><RANKING place="5" resultid="3520"/><RANKING place="6" resultid="3522"/><RANKING place="9" resultid="3528"/><RANKING place="3" resultid="3533"/><RANKING place="2" resultid="3540"/><RANKING place="4" resultid="3542"/><RANKING place="1" resultid="3555"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="400009" agemax="16" agemin="16" gender="M" name="Jahrgang 2009"><RANKINGS><RANKING place="17" resultid="3495"/><RANKING place="12" resultid="3500"/><RANKING place="-1" resultid="3505"/><RANKING place="15" resultid="3507"/><RANKING place="14" resultid="3513"/><RANKING place="18" resultid="3517"/><RANKING place="6" resultid="3524"/><RANKING place="13" resultid="3525"/><RANKING place="8" resultid="3526"/><RANKING place="16" resultid="3529"/><RANKING place="2" resultid="3531"/><RANKING place="9" resultid="3535"/><RANKING place="11" resultid="3536"/><RANKING place="4" resultid="3541"/><RANKING place="1" resultid="3546"/><RANKING place="7" resultid="3547"/><RANKING place="3" resultid="3548"/><RANKING place="5" resultid="3549"/><RANKING place="10" resultid="3557"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="400010" agemax="17" agemin="17" gender="M" name="Jahrgang 2008"><RANKINGS><RANKING place="4" resultid="3442"/><RANKING place="6" resultid="3498"/><RANKING place="-1" resultid="3523"/><RANKING place="5" resultid="3527"/><RANKING place="2" resultid="3538"/><RANKING place="3" resultid="3551"/><RANKING place="1" resultid="3553"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="400011" agemax="-1" agemin="18" gender="M" name="Jahrgang 2007 und älter"><RANKINGS><RANKING place="15" resultid="3503"/><RANKING place="13" resultid="3511"/><RANKING place="14" resultid="3516"/><RANKING place="10" resultid="3519"/><RANKING place="-1" resultid="3521"/><RANKING place="6" resultid="3532"/><RANKING place="9" resultid="3534"/><RANKING place="8" resultid="3539"/><RANKING place="7" resultid="3544"/><RANKING place="11" resultid="3545"/><RANKING place="5" resultid="3550"/><RANKING place="4" resultid="3552"/><RANKING place="3" resultid="3554"/><RANKING place="1" resultid="3556"/><RANKING place="12" resultid="3558"/><RANKING place="2" resultid="3559"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="451" number="1" order="1" status="OFFICIAL"/><HEAT heatid="452" number="2" order="2" status="OFFICIAL"/><HEAT heatid="453" number="3" order="3" status="OFFICIAL"/><HEAT heatid="454" number="4" order="4" status="OFFICIAL"/><HEAT heatid="455" number="5" order="5" status="OFFICIAL"/><HEAT heatid="456" number="6" order="6" status="OFFICIAL"/><HEAT heatid="457" number="7" order="7" status="OFFICIAL"/><HEAT heatid="458" number="8" order="8" status="OFFICIAL"/><HEAT heatid="459" number="9" order="9" status="OFFICIAL"/><HEAT heatid="460" number="10" order="10" status="OFFICIAL"/><HEAT heatid="461" number="11" order="11" status="OFFICIAL"/><HEAT heatid="462" number="12" order="12" status="OFFICIAL"/><HEAT heatid="463" number="13" order="13" status="OFFICIAL"/><HEAT heatid="464" number="14" order="14" status="OFFICIAL"/><HEAT heatid="465" number="15" order="15" status="OFFICIAL"/><HEAT heatid="466" number="16" order="16" status="OFFICIAL"/><HEAT heatid="467" number="17" order="17" status="OFFICIAL"/><HEAT heatid="468" number="18" order="18" status="OFFICIAL"/><HEAT heatid="469" number="19" order="19" status="OFFICIAL"/><HEAT heatid="470" number="20" order="20" status="OFFICIAL"/><HEAT heatid="471" number="21" order="21" status="OFFICIAL"/><HEAT heatid="472" number="22" order="22" status="OFFICIAL"/><HEAT heatid="473" number="23" order="23" status="OFFICIAL"/><HEAT heatid="474" number="24" order="24" status="OFFICIAL"/><HEAT heatid="475" number="25" order="25" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT><EVENT eventid="41" gender="F" number="41" order="41" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="700"/><SWIMSTYLE distance="400" name="400m Lagen Frauen" relaycount="1" stroke="MEDLEY"/><AGEGROUPS><AGEGROUP agegroupid="410001" agemax="11" agemin="11" gender="F" name="Jahrgang 2014"><RANKINGS><RANKING place="1" resultid="3562"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="410002" agemax="12" agemin="12" gender="F" name="Jahrgang 2013"><RANKINGS><RANKING place="2" resultid="3560"/><RANKING place="1" resultid="3563"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="410003" agemax="13" agemin="13" gender="F" name="Jahrgang 2012"><RANKINGS><RANKING place="1" resultid="3567"/><RANKING place="2" resultid="3569"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="410004" agemax="14" agemin="14" gender="F" name="Jahrgang 2011"><RANKINGS><RANKING place="2" resultid="3565"/><RANKING place="3" resultid="3566"/><RANKING place="1" resultid="3570"/><RANKING place="4" resultid="3577"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="410005" agemax="15" agemin="15" gender="F" name="Jahrgang 2010"><RANKINGS><RANKING place="3" resultid="3561"/><RANKING place="2" resultid="3564"/><RANKING place="1" resultid="3575"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="410006" agemax="16" agemin="16" gender="F" name="Jahrgang 2009"><RANKINGS><RANKING place="1" resultid="3571"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="410007" agemax="17" agemin="17" gender="F" name="Jahrgang 2008"><RANKINGS><RANKING place="1" resultid="3572"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="410008" agemax="-1" agemin="18" gender="F" name="Jahrgang 2007 und älter"><RANKINGS><RANKING place="3" resultid="3568"/><RANKING place="1" resultid="3573"/><RANKING place="2" resultid="3574"/><RANKING place="4" resultid="3576"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="476" number="1" order="1" status="OFFICIAL"/><HEAT heatid="477" number="2" order="2" status="OFFICIAL"/><HEAT heatid="478" number="3" order="3" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT><EVENT eventid="42" gender="M" number="42" order="42" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="ATHLETE" value="700"/><SWIMSTYLE distance="400" name="400m Lagen Männer" relaycount="1" stroke="MEDLEY"/><AGEGROUPS><AGEGROUP agegroupid="420001" agemax="11" agemin="11" gender="M" name="Jahrgang 2014"><RANKINGS/></AGEGROUP><AGEGROUP agegroupid="420002" agemax="12" agemin="12" gender="M" name="Jahrgang 2013"><RANKINGS><RANKING place="1" resultid="3584"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="420003" agemax="13" agemin="13" gender="M" name="Jahrgang 2012"><RANKINGS><RANKING place="-1" resultid="3578"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="420004" agemax="14" agemin="14" gender="M" name="Jahrgang 2011"><RANKINGS><RANKING place="2" resultid="3581"/><RANKING place="-1" resultid="3586"/><RANKING place="3" resultid="3590"/><RANKING place="1" resultid="3591"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="420005" agemax="15" agemin="15" gender="M" name="Jahrgang 2010"><RANKINGS><RANKING place="6" resultid="3580"/><RANKING place="4" resultid="3585"/><RANKING place="3" resultid="3587"/><RANKING place="5" resultid="3588"/><RANKING place="7" resultid="3589"/><RANKING place="2" resultid="3593"/><RANKING place="1" resultid="3596"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="420006" agemax="16" agemin="16" gender="M" name="Jahrgang 2009"><RANKINGS><RANKING place="1" resultid="3579"/><RANKING place="4" resultid="3582"/><RANKING place="3" resultid="3583"/><RANKING place="2" resultid="3592"/></RANKINGS></AGEGROUP><AGEGROUP agegroupid="420007" agemax="17" agemin="17" gender="M" name="Jahrgang 2008"><RANKINGS/></AGEGROUP><AGEGROUP agegroupid="420008" agemax="-1" agemin="18" gender="M" name="Jahrgang 2007 und älter"><RANKINGS><RANKING place="1" resultid="3594"/><RANKING place="2" resultid="3595"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="479" number="1" order="1" status="OFFICIAL"/><HEAT heatid="480" number="2" order="2" status="OFFICIAL"/><HEAT heatid="481" number="3" order="3" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT><EVENT eventid="43" gender="F" number="43" order="43" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="RELAY" value="2500"/><SWIMSTYLE distance="200" name="4x200m Freistil Frauen" relaycount="4" stroke="FREE"/><AGEGROUPS><AGEGROUP agegroupid="430001" agemax="-1" agemin="9" gender="F" name="Jahrgang 2016 und älter"><RANKINGS><RANKING place="1" resultid="3597"/><RANKING place="2" resultid="3598"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="482" number="1" order="1" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT><EVENT eventid="44" gender="M" number="44" order="44" round="TIM" timing="AUTOMATIC"><FEE currency="EUR" type="RELAY" value="2500"/><SWIMSTYLE distance="200" name="4x200m Freistil Männer" relaycount="4" stroke="FREE"/><AGEGROUPS><AGEGROUP agegroupid="440001" agemax="-1" agemin="9" gender="M" name="Jahrgang 2016 und älter"><RANKINGS><RANKING place="1" resultid="3599"/></RANKINGS></AGEGROUP></AGEGROUPS><HEATS><HEAT heatid="483" number="1" order="1" status="OFFICIAL"/></HEATS><TIMESTANDARDREFS/></EVENT></EVENTS></SESSION></SESSIONS><CLUBS><CLUB code="4392" name="TB Erlangen" nation="GER" region="02" shortname="TBErl" type="CLUB"><CONTACT city="Erlangen" email="meldungen.schwimmen@tb-erlangen.de" name="Zebelein, Christian" phone="+49 176 32619612" street="Nägelsbachstr. 27" zip="91052"/><OFFICIALS/><ATHLETES><ATHLETE athleteid="1" birthdate="2013-01-01" firstname="Helena" gender="F" lastname="Kurtz" license="504316"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="1" lane="3" resultid="1" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="9" heatid="102" lane="4" resultid="766" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="27" heatid="253" lane="8" resultid="1875" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="31" heatid="327" lane="3" resultid="2430" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="2" birthdate="2015-01-01" firstname="Shriya" gender="F" lastname="Badrinarayanan" license="504318"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="1" lane="4" points="57" resultid="2" swimtime="00:01:16.08"><SPLITS/></RESULT><RESULT eventid="9" heatid="102" lane="6" points="54" resultid="768" swimtime="00:01:02.40"><SPLITS/></RESULT><RESULT eventid="27" heatid="252" lane="6" points="60" resultid="1866" swimtime="00:01:08.67"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="3" birthdate="2014-01-01" firstname="Elena" gender="F" lastname="Vojtisek" license="504302"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="1" lane="5" points="182" resultid="3" swimtime="00:00:51.68"><SPLITS/></RESULT><RESULT eventid="9" heatid="102" lane="2" points="164" resultid="764" swimtime="00:00:43.21"><SPLITS/></RESULT><RESULT eventid="23" heatid="240" lane="5" resultid="1792" swimtime="00:00:58.72"><SPLITS/></RESULT><RESULT eventid="27" heatid="252" lane="5" points="143" resultid="1865" swimtime="00:00:51.53"><SPLITS/></RESULT><RESULT eventid="39" heatid="420" lane="3" points="130" resultid="3127" swimtime="00:01:41.89"><SPLITS><SPLIT distance="50" swimtime="00:00:45.29"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="4" birthdate="2012-01-01" firstname="Shin" gender="F" lastname="Lee" license="504323"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="1" lane="6" points="243" resultid="4" swimtime="00:00:46.89"><SPLITS/></RESULT><RESULT eventid="9" heatid="102" lane="3" points="155" resultid="765" swimtime="00:00:44.03"><SPLITS/></RESULT><RESULT eventid="27" heatid="252" lane="7" points="129" resultid="1867" swimtime="00:00:53.31"><SPLITS/></RESULT><RESULT eventid="31" heatid="327" lane="7" points="241" resultid="2434" swimtime="00:01:43.04"><SPLITS><SPLIT distance="50" swimtime="00:00:49.35"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="5" birthdate="2011-01-01" firstname="Leonie" gender="F" lastname="Balling" license="504304"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="2" lane="1" points="275" resultid="5" swimtime="00:00:45.01"><SPLITS/></RESULT><RESULT eventid="9" heatid="103" lane="1" points="293" resultid="769" swimtime="00:00:35.61"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="6" birthdate="2013-01-01" firstname="Kavya" gender="F" lastname="Jeyavelan" license="504322"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="2" lane="2" points="143" resultid="6" swimtime="00:00:55.99"><SPLITS/></RESULT><RESULT eventid="9" heatid="103" lane="8" points="110" resultid="776" swimtime="00:00:49.32"><SPLITS/></RESULT><RESULT eventid="27" heatid="252" lane="2" points="91" resultid="1862" swimtime="00:00:59.90"><SPLITS/></RESULT><RESULT eventid="31" heatid="326" lane="3" points="117" resultid="2426" swimtime="00:02:10.78"><SPLITS><SPLIT distance="50" swimtime="00:01:03.42"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="7" birthdate="2017-01-01" firstname="Bella" gender="F" lastname="Buchert" license="504243"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="2" lane="3" points="97" resultid="7" swimtime="00:01:03.67"><SPLITS/></RESULT><RESULT eventid="9" heatid="103" lane="2" points="32" resultid="770" swimtime="00:01:14.21"><SPLITS/></RESULT><RESULT eventid="27" heatid="253" lane="1" points="59" resultid="1868" swimtime="00:01:09.10"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="8" birthdate="2017-01-01" firstname="Paula" gender="F" lastname="Moosmeier" license="504242"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="2" lane="4" points="93" resultid="8" swimtime="00:01:04.56"><SPLITS/></RESULT><RESULT eventid="27" heatid="253" lane="7" points="55" resultid="1874" swimtime="00:01:10.66"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="10" birthdate="2014-01-01" firstname="Laura" gender="F" lastname="De Andrews" license="504319"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="2" lane="6" points="90" resultid="10" swimtime="00:01:05.31"><SPLITS/></RESULT><RESULT eventid="9" heatid="102" lane="5" points="88" resultid="767" swimtime="00:00:53.02"><SPLITS/></RESULT><RESULT eventid="25" heatid="246" lane="3" resultid="1828" swimtime="00:01:13.84"><SPLITS/></RESULT><RESULT eventid="27" heatid="252" lane="3" points="85" resultid="1863" swimtime="00:01:01.17"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="11" birthdate="2015-01-01" firstname="Diya" gender="F" lastname="Jeyavelan" license="504321"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="2" lane="7" points="88" resultid="11" swimtime="00:01:05.64"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="12" birthdate="2015-01-01" firstname="Melina" gender="F" lastname="Madhan" license="504324"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="2" lane="8" points="77" resultid="12" swimtime="00:01:08.68"><SPLITS/></RESULT><RESULT eventid="27" heatid="252" lane="4" points="46" resultid="1864" swimtime="00:01:14.89"><SPLITS/></RESULT><RESULT eventid="31" heatid="326" lane="5" points="90" resultid="2428" swimtime="00:02:22.84"><SPLITS><SPLIT distance="50" swimtime="00:01:04.52"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="14" birthdate="2013-01-01" firstname="Minou" gender="F" lastname="Köhl" license="504244"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="3" lane="2" resultid="14" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="9" heatid="103" lane="3" resultid="771" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="27" heatid="253" lane="5" resultid="1872" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="17" birthdate="2013-01-01" firstname="Lotta" gender="F" lastname="Blum" license="470677"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="3" lane="5" points="125" resultid="17" swimtime="00:00:58.46"><SPLITS/></RESULT><RESULT eventid="9" heatid="104" lane="2" points="118" resultid="778" swimtime="00:00:48.17"><SPLITS/></RESULT><RESULT eventid="27" heatid="254" lane="1" points="115" resultid="1876" swimtime="00:00:55.39"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="18" birthdate="2014-01-01" firstname="Moira" gender="F" lastname="Baxter" license="470850"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="3" lane="6" points="141" resultid="18" swimtime="00:00:56.17"><SPLITS/></RESULT><RESULT eventid="25" heatid="246" lane="5" resultid="1830" swimtime="00:01:02.99"><SPLITS/></RESULT><RESULT eventid="31" heatid="326" lane="4" points="120" resultid="2427" swimtime="00:02:09.91"><SPLITS><SPLIT distance="50" swimtime="00:01:01.97"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="19" birthdate="2016-01-01" firstname="Astrid" gender="F" lastname="van de Stadt" license="498610"><HANDICAP/><ENTRIES/><RESULTS><RESULT comment="09:13 Der Zielanschlag erfolgte nicht mit beiden Händen gleichzeitig" eventid="1" heatid="3" lane="7" resultid="19" status="DSQ" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="9" heatid="103" lane="6" points="57" resultid="774" swimtime="00:01:01.44"><SPLITS/></RESULT><RESULT eventid="27" heatid="253" lane="3" points="80" resultid="1870" swimtime="00:01:02.41"><SPLITS/></RESULT><RESULT eventid="39" heatid="421" lane="8" points="54" resultid="3138" swimtime="00:02:16.46"><SPLITS><SPLIT distance="50" swimtime="00:01:06.37"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="22" birthdate="2016-01-01" firstname="Maja" gender="F" lastname="Hagen" license="491452"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="4" lane="2" points="142" resultid="22" swimtime="00:00:56.07"><SPLITS/></RESULT><RESULT eventid="9" heatid="109" lane="4" points="191" resultid="820" swimtime="00:00:41.07"><SPLITS/></RESULT><RESULT eventid="13" heatid="194" lane="5" points="164" resultid="1468" swimtime="00:01:44.90"><SPLITS><SPLIT distance="50" swimtime="00:00:53.58"/></SPLITS></RESULT><RESULT eventid="27" heatid="256" lane="6" points="186" resultid="1897" swimtime="00:00:47.19"><SPLITS/></RESULT><RESULT eventid="29" heatid="290" lane="5" points="164" resultid="2155" swimtime="00:03:26.21"><SPLITS><SPLIT distance="50" swimtime="00:00:46.87"/><SPLIT distance="100" swimtime="00:01:41.21"/><SPLIT distance="150" swimtime="00:02:36.34"/></SPLITS></RESULT><RESULT eventid="35" heatid="364" lane="1" points="104" resultid="2703" swimtime="00:00:51.84"><SPLITS/></RESULT><RESULT eventid="39" heatid="426" lane="3" points="165" resultid="3172" swimtime="00:01:34.22"><SPLITS><SPLIT distance="50" swimtime="00:00:45.82"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="24" birthdate="2016-01-01" firstname="Elena" gender="F" lastname="Barozzi" license="495062"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="4" lane="4" points="104" resultid="24" swimtime="00:01:02.19"><SPLITS/></RESULT><RESULT eventid="9" heatid="103" lane="4" points="100" resultid="772" swimtime="00:00:50.87"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="25" birthdate="2017-01-01" firstname="Isabelle" gender="F" lastname="Möbus" license="490446"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="4" lane="5" points="111" resultid="25" swimtime="00:01:00.90"><SPLITS/></RESULT><RESULT eventid="9" heatid="104" lane="3" points="96" resultid="779" swimtime="00:00:51.58"><SPLITS/></RESULT><RESULT eventid="13" heatid="192" lane="6" points="81" resultid="1453" swimtime="00:02:12.54"><SPLITS><SPLIT distance="50" swimtime="00:01:01.30"/></SPLITS></RESULT><RESULT eventid="27" heatid="254" lane="8" points="96" resultid="1883" swimtime="00:00:58.89"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="26" birthdate="2016-01-01" firstname="Antonina" gender="F" lastname="Lukina" license="495021"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="4" lane="6" points="104" resultid="26" swimtime="00:01:02.26"><SPLITS/></RESULT><RESULT comment="14:10 Start vor dem Startsignal" eventid="9" heatid="105" lane="8" resultid="792" status="DSQ" swimtime="NT"><SPLITS/></RESULT><RESULT comment="16:52 Start vor dem Startsignal" eventid="13" heatid="191" lane="3" resultid="1442" status="DSQ" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="27" heatid="255" lane="8" points="120" resultid="1891" swimtime="00:00:54.59"><SPLITS/></RESULT><RESULT eventid="39" heatid="422" lane="1" points="111" resultid="3139" swimtime="00:01:47.54"><SPLITS><SPLIT distance="50" swimtime="00:00:50.70"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="29" birthdate="2015-01-01" firstname="Alexandra" gender="F" lastname="Brussilowski" license="479245"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="5" lane="1" points="120" resultid="29" swimtime="00:00:59.29"><SPLITS/></RESULT><RESULT comment="14:09 Start vor dem Startsignal" eventid="9" heatid="106" lane="8" resultid="800" status="DSQ" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="13" heatid="191" lane="7" points="115" resultid="1446" swimtime="00:01:58.02"><SPLITS><SPLIT distance="50" swimtime="00:00:58.70"/></SPLITS></RESULT><RESULT eventid="27" heatid="256" lane="8" points="97" resultid="1899" swimtime="00:00:58.64"><SPLITS/></RESULT><RESULT eventid="39" heatid="422" lane="6" points="112" resultid="3144" swimtime="00:01:47.10"><SPLITS><SPLIT distance="50" swimtime="00:00:50.81"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="36" birthdate="2017-01-01" firstname="Emma" gender="F" lastname="Zhuang" license="499826"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="5" lane="8" points="99" resultid="36" swimtime="00:01:03.17"><SPLITS/></RESULT><RESULT eventid="9" heatid="104" lane="7" points="133" resultid="783" swimtime="00:00:46.37"><SPLITS/></RESULT><RESULT eventid="13" heatid="192" lane="3" points="130" resultid="1450" swimtime="00:01:53.12"><SPLITS><SPLIT distance="50" swimtime="00:00:54.36"/></SPLITS></RESULT><RESULT eventid="27" heatid="254" lane="5" points="109" resultid="1880" swimtime="00:00:56.33"><SPLITS/></RESULT><RESULT eventid="39" heatid="421" lane="1" points="111" resultid="3131" swimtime="00:01:47.32"><SPLITS><SPLIT distance="50" swimtime="00:00:49.80"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="45" birthdate="2016-01-01" firstname="Halina" gender="F" lastname="Kojro" license="485126"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="7" lane="1" points="133" resultid="45" swimtime="00:00:57.26"><SPLITS/></RESULT><RESULT eventid="9" heatid="108" lane="4" points="199" resultid="812" swimtime="00:00:40.54"><SPLITS/></RESULT><RESULT eventid="13" heatid="195" lane="6" points="216" resultid="1477" swimtime="00:01:35.61"><SPLITS><SPLIT distance="50" swimtime="00:00:46.63"/></SPLITS></RESULT><RESULT eventid="27" heatid="260" lane="7" points="200" resultid="1930" swimtime="00:00:46.07"><SPLITS/></RESULT><RESULT eventid="35" heatid="365" lane="3" points="154" resultid="2713" swimtime="00:00:45.56"><SPLITS/></RESULT><RESULT eventid="37" heatid="403" lane="6" points="208" resultid="3004" swimtime="00:03:28.09"><SPLITS><SPLIT distance="50" swimtime="00:00:49.51"/><SPLIT distance="100" swimtime="00:01:44.17"/><SPLIT distance="150" swimtime="00:02:37.84"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="49" birthdate="2015-01-01" firstname="Josefine Mia" gender="F" lastname="Felderer" license="495022"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="7" lane="5" points="171" resultid="49" swimtime="00:00:52.70"><SPLITS/></RESULT><RESULT eventid="9" heatid="106" lane="3" points="123" resultid="795" swimtime="00:00:47.57"><SPLITS/></RESULT><RESULT eventid="27" heatid="256" lane="7" points="160" resultid="1898" swimtime="00:00:49.64"><SPLITS/></RESULT><RESULT eventid="31" heatid="329" lane="2" points="139" resultid="2444" swimtime="00:02:03.62"><SPLITS><SPLIT distance="50" swimtime="00:00:59.67"/></SPLITS></RESULT><RESULT eventid="39" heatid="422" lane="8" points="115" resultid="3146" swimtime="00:01:46.10"><SPLITS><SPLIT distance="50" swimtime="00:00:51.65"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="52" birthdate="2015-01-01" firstname="Selma Ruth" gender="F" lastname="Jannack" license="499857"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="7" lane="8" points="112" resultid="52" swimtime="00:01:00.69"><SPLITS/></RESULT><RESULT eventid="9" heatid="107" lane="1" points="129" resultid="801" swimtime="00:00:46.77"><SPLITS/></RESULT><RESULT eventid="13" heatid="192" lane="5" resultid="1452" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="27" heatid="255" lane="3" points="150" resultid="1886" swimtime="00:00:50.71"><SPLITS/></RESULT><RESULT comment="10:00 Die Sportlerin hat nicht die vollständige Wettkampfstrecke absolviert" eventid="29" heatid="288" lane="6" resultid="2142" status="DSQ" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="39" heatid="421" lane="5" points="123" resultid="3135" swimtime="00:01:43.91"><SPLITS><SPLIT distance="50" swimtime="00:00:47.84"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="57" birthdate="2016-01-01" firstname="Viktoria" gender="F" lastname="Nagy" license="488904"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="8" lane="5" points="208" resultid="57" swimtime="00:00:49.40"><SPLITS/></RESULT><RESULT eventid="9" heatid="111" lane="1" points="222" resultid="833" swimtime="00:00:39.07"><SPLITS/></RESULT><RESULT eventid="13" heatid="196" lane="8" points="178" resultid="1487" swimtime="00:01:42.08"><SPLITS><SPLIT distance="50" swimtime="00:00:51.33"/></SPLITS></RESULT><RESULT eventid="29" heatid="293" lane="8" points="235" resultid="2181" swimtime="00:03:03.02"><SPLITS><SPLIT distance="50" swimtime="00:00:42.08"/><SPLIT distance="100" swimtime="00:01:28.92"/><SPLIT distance="150" swimtime="00:02:18.91"/></SPLITS></RESULT><RESULT eventid="31" heatid="332" lane="8" points="198" resultid="2474" swimtime="00:01:49.98"><SPLITS><SPLIT distance="50" swimtime="00:00:53.47"/></SPLITS></RESULT><RESULT eventid="37" heatid="403" lane="3" points="193" resultid="3001" swimtime="00:03:33.15"><SPLITS><SPLIT distance="50" swimtime="00:00:49.73"/><SPLIT distance="100" swimtime="00:01:45.18"/><SPLIT distance="150" swimtime="00:02:40.31"/></SPLITS></RESULT><RESULT eventid="39" heatid="427" lane="2" points="192" resultid="3179" swimtime="00:01:29.62"><SPLITS><SPLIT distance="50" swimtime="00:00:43.06"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="62" birthdate="2015-01-01" firstname="Valentina" gender="F" lastname="Plenkers" license="479303"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="9" lane="2" points="119" resultid="62" swimtime="00:00:59.45"><SPLITS/></RESULT><RESULT eventid="9" heatid="107" lane="3" points="173" resultid="803" swimtime="00:00:42.40"><SPLITS/></RESULT><RESULT eventid="27" heatid="255" lane="6" points="139" resultid="1889" swimtime="00:00:52.02"><SPLITS/></RESULT><RESULT eventid="29" heatid="289" lane="4" points="151" resultid="2146" swimtime="00:03:32.15"><SPLITS><SPLIT distance="50" swimtime="00:00:49.14"/><SPLIT distance="100" swimtime="00:01:45.30"/><SPLIT distance="150" swimtime="00:02:42.46"/></SPLITS></RESULT><RESULT eventid="35" heatid="364" lane="7" points="47" resultid="2709" swimtime="00:01:07.59"><SPLITS/></RESULT><RESULT eventid="39" heatid="425" lane="6" points="144" resultid="3167" swimtime="00:01:38.53"><SPLITS><SPLIT distance="50" swimtime="00:00:47.26"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="73" birthdate="2013-01-01" firstname="Thuy An" gender="F" lastname="Nguyen" license="460255"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="10" lane="5" points="254" resultid="73" swimtime="00:00:46.23"><SPLITS/></RESULT><RESULT eventid="9" heatid="105" lane="7" points="160" resultid="791" swimtime="00:00:43.58"><SPLITS/></RESULT><RESULT eventid="25" heatid="247" lane="2" resultid="1831" swimtime="00:00:54.89"><SPLITS/></RESULT><RESULT eventid="31" heatid="331" lane="5" points="266" resultid="2463" swimtime="00:01:39.62"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="78" birthdate="2013-01-01" firstname="Katja" gender="F" lastname="Khodyachykh" license="479063"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="11" lane="2" points="195" resultid="78" swimtime="00:00:50.46"><SPLITS/></RESULT><RESULT eventid="9" heatid="110" lane="3" points="223" resultid="827" swimtime="00:00:39.01"><SPLITS/></RESULT><RESULT eventid="25" heatid="246" lane="4" resultid="1829" swimtime="00:01:01.44"><SPLITS/></RESULT><RESULT eventid="27" heatid="258" lane="5" points="147" resultid="1912" swimtime="00:00:51.01"><SPLITS/></RESULT><RESULT eventid="31" heatid="333" lane="5" points="191" resultid="2479" swimtime="00:01:51.26"><SPLITS><SPLIT distance="50" swimtime="00:00:51.27"/></SPLITS></RESULT><RESULT eventid="39" heatid="421" lane="3" points="154" resultid="3133" swimtime="00:01:36.43"><SPLITS><SPLIT distance="50" swimtime="00:00:46.01"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="187" birthdate="2013-01-01" firstname="Emil" gender="M" lastname="Biondic" license="504303"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="25" lane="3" points="114" resultid="187" swimtime="00:00:53.43"><SPLITS/></RESULT><RESULT eventid="10" heatid="133" lane="2" points="142" resultid="1000" swimtime="00:00:40.02"><SPLITS/></RESULT><RESULT eventid="26" heatid="250" lane="5" resultid="1855" swimtime="00:01:00.80"><SPLITS/></RESULT><RESULT eventid="32" heatid="345" lane="3" points="125" resultid="2571" swimtime="00:01:53.47"><SPLITS><SPLIT distance="50" swimtime="00:00:53.95"/></SPLITS></RESULT><RESULT eventid="40" heatid="451" lane="3" points="118" resultid="3368" swimtime="00:01:35.51"><SPLITS><SPLIT distance="50" swimtime="00:00:44.70"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="188" birthdate="2017-01-01" firstname="Torge" gender="M" lastname="Rießland" license="504132"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="25" lane="4" points="53" resultid="188" swimtime="00:01:08.85"><SPLITS/></RESULT><RESULT eventid="10" heatid="133" lane="6" points="30" resultid="1004" swimtime="00:01:07.22"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="189" birthdate="2017-01-01" firstname="Louis" gender="M" lastname="Lambertus" license="504589"><HANDICAP/><ENTRIES/><RESULTS><RESULT comment="09:37 Start vor dem Startsignal" eventid="2" heatid="25" lane="5" resultid="189" status="DSQ" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="190" birthdate="2016-01-01" firstname="Tom" gender="M" lastname="Reuling" license="504133"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="26" lane="1" points="60" resultid="190" swimtime="00:01:06.17"><SPLITS/></RESULT><RESULT eventid="10" heatid="133" lane="3" points="44" resultid="1001" swimtime="00:00:59.07"><SPLITS/></RESULT><RESULT eventid="28" heatid="274" lane="1" points="57" resultid="2031" swimtime="00:01:01.49"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="191" birthdate="2016-01-01" firstname="Anton" gender="M" lastname="Träbing" license="504817"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="26" lane="2" resultid="191" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="192" birthdate="2016-01-01" firstname="Max" gender="M" lastname="Splihal" license="495067"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="26" lane="3" points="58" resultid="192" swimtime="00:01:07.02"><SPLITS/></RESULT><RESULT eventid="10" heatid="134" lane="8" points="53" resultid="1012" swimtime="00:00:55.58"><SPLITS/></RESULT><RESULT eventid="14" heatid="210" lane="7" points="78" resultid="1596" swimtime="00:02:00.30"><SPLITS><SPLIT distance="50" swimtime="00:00:57.20"/></SPLITS></RESULT><RESULT eventid="28" heatid="274" lane="2" points="66" resultid="2032" swimtime="00:00:58.64"><SPLITS/></RESULT><RESULT eventid="40" heatid="452" lane="1" points="67" resultid="3374" swimtime="00:01:55.25"><SPLITS><SPLIT distance="50" swimtime="00:00:56.82"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="196" birthdate="2016-01-01" firstname="Laurens" gender="M" lastname="Lambertus" license="504588"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="26" lane="7" points="67" resultid="196" swimtime="00:01:03.69"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="197" birthdate="2016-01-01" firstname="Moritz" gender="M" lastname="Köhl" license="504245"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="26" lane="8" points="69" resultid="197" swimtime="00:01:03.20"><SPLITS/></RESULT><RESULT eventid="10" heatid="133" lane="5" points="42" resultid="1003" swimtime="00:01:00.06"><SPLITS/></RESULT><RESULT eventid="28" heatid="274" lane="8" points="42" resultid="2038" swimtime="00:01:07.85"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="200" birthdate="2015-01-01" firstname="Eric" gender="M" lastname="Rosu" license="494783"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="27" lane="3" points="114" resultid="200" swimtime="00:00:53.40"><SPLITS/></RESULT><RESULT eventid="10" heatid="134" lane="6" points="87" resultid="1010" swimtime="00:00:47.14"><SPLITS/></RESULT><RESULT eventid="14" heatid="210" lane="3" points="102" resultid="1592" swimtime="00:01:50.08"><SPLITS><SPLIT distance="50" swimtime="00:00:53.15"/></SPLITS></RESULT><RESULT eventid="28" heatid="275" lane="6" points="114" resultid="2044" swimtime="00:00:48.82"><SPLITS/></RESULT><RESULT eventid="30" heatid="309" lane="6" points="72" resultid="2301" swimtime="00:04:04.63"><SPLITS><SPLIT distance="50" swimtime="00:00:53.85"/><SPLIT distance="100" swimtime="00:01:59.01"/><SPLIT distance="150" swimtime="00:03:05.20"/></SPLITS></RESULT><RESULT eventid="40" heatid="452" lane="7" points="85" resultid="3380" swimtime="00:01:46.45"><SPLITS><SPLIT distance="50" swimtime="00:00:49.29"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="202" birthdate="2015-01-01" firstname="Eric" gender="M" lastname="Lütcke" license="489959"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="27" lane="5" points="83" resultid="202" swimtime="00:00:59.40"><SPLITS/></RESULT><RESULT eventid="10" heatid="134" lane="5" points="88" resultid="1009" swimtime="00:00:46.98"><SPLITS/></RESULT><RESULT eventid="28" heatid="274" lane="6" points="77" resultid="2036" swimtime="00:00:55.63"><SPLITS/></RESULT><RESULT eventid="30" heatid="309" lane="7" points="69" resultid="2302" swimtime="00:04:07.63"><SPLITS><SPLIT distance="50" swimtime="00:00:52.38"/><SPLIT distance="100" swimtime="00:02:00.75"/><SPLIT distance="150" swimtime="00:03:05.73"/></SPLITS></RESULT><RESULT eventid="40" heatid="453" lane="7" points="77" resultid="3388" swimtime="00:01:49.85"><SPLITS><SPLIT distance="50" swimtime="00:00:51.27"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="203" birthdate="2016-01-01" firstname="Haobin" gender="M" lastname="Sun" license="485142"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="27" lane="7" points="118" resultid="203" swimtime="00:00:52.78"><SPLITS/></RESULT><RESULT eventid="10" heatid="133" lane="4" points="90" resultid="1002" swimtime="00:00:46.52"><SPLITS/></RESULT><RESULT eventid="28" heatid="274" lane="5" points="92" resultid="2035" swimtime="00:00:52.51"><SPLITS/></RESULT><RESULT eventid="40" heatid="452" lane="3" points="80" resultid="3376" swimtime="00:01:48.73"><SPLITS><SPLIT distance="50" swimtime="00:00:52.54"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="209" birthdate="2015-01-01" firstname="Noah Nikolas" gender="M" lastname="Wicklein" license="498832"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="28" lane="5" points="95" resultid="209" swimtime="00:00:56.87"><SPLITS/></RESULT><RESULT eventid="10" heatid="135" lane="5" points="109" resultid="1017" swimtime="00:00:43.69"><SPLITS/></RESULT><RESULT eventid="14" heatid="210" lane="4" points="106" resultid="1593" swimtime="00:01:48.71"><SPLITS><SPLIT distance="50" swimtime="00:00:52.69"/></SPLITS></RESULT><RESULT eventid="28" heatid="274" lane="4" points="109" resultid="2034" swimtime="00:00:49.58"><SPLITS/></RESULT><RESULT eventid="40" heatid="452" lane="5" points="102" resultid="3378" swimtime="00:01:40.04"><SPLITS><SPLIT distance="50" swimtime="00:00:45.49"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="215" birthdate="2014-01-01" firstname="Valentin" gender="M" lastname="Gopych" license="475139"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="29" lane="3" points="118" resultid="215" swimtime="00:00:52.80"><SPLITS/></RESULT><RESULT eventid="10" heatid="134" lane="7" points="96" resultid="1011" swimtime="00:00:45.66"><SPLITS/></RESULT><RESULT eventid="22" heatid="239" lane="2" resultid="1785" swimtime="00:01:18.78"><SPLITS/></RESULT><RESULT eventid="28" heatid="275" lane="8" points="76" resultid="2046" swimtime="00:00:55.91"><SPLITS/></RESULT><RESULT eventid="32" heatid="346" lane="8" points="109" resultid="2581" swimtime="00:01:58.78"><SPLITS><SPLIT distance="50" swimtime="00:00:54.27"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="227" birthdate="2015-01-01" firstname="Emanuel" gender="M" lastname="Hauer" license="488589"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="30" lane="7" points="159" resultid="227" swimtime="00:00:47.85"><SPLITS/></RESULT><RESULT eventid="10" heatid="136" lane="1" points="121" resultid="1021" swimtime="00:00:42.24"><SPLITS/></RESULT><RESULT eventid="28" heatid="275" lane="2" points="107" resultid="2040" swimtime="00:00:49.81"><SPLITS/></RESULT><RESULT eventid="30" heatid="310" lane="3" points="95" resultid="2306" swimtime="00:03:43.03"><SPLITS><SPLIT distance="50" swimtime="00:00:44.85"/><SPLIT distance="100" swimtime="00:01:43.51"/><SPLIT distance="150" swimtime="00:02:44.87"/></SPLITS></RESULT><RESULT eventid="36" heatid="385" lane="1" points="66" resultid="2863" swimtime="00:00:54.84"><SPLITS/></RESULT><RESULT eventid="40" heatid="453" lane="3" points="112" resultid="3384" swimtime="00:01:37.05"><SPLITS><SPLIT distance="50" swimtime="00:00:44.70"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="510" birthdate="2015-01-01" firstname="Aaron" gender="M" lastname="Hoffmann" license="487806"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="8" heatid="93" lane="4" points="172" resultid="700" swimtime="00:03:46.30"><SPLITS><SPLIT distance="50" swimtime="00:00:52.31"/><SPLIT distance="100" swimtime="00:01:50.56"/><SPLIT distance="150" swimtime="00:02:48.86"/></SPLITS></RESULT><RESULT eventid="10" heatid="135" lane="6" points="119" resultid="1018" swimtime="00:00:42.50"><SPLITS/></RESULT><RESULT eventid="14" heatid="214" lane="1" points="174" resultid="1621" swimtime="00:01:32.27"><SPLITS><SPLIT distance="50" swimtime="00:00:45.83"/></SPLITS></RESULT><RESULT eventid="28" heatid="277" lane="6" points="148" resultid="2058" swimtime="00:00:44.74"><SPLITS/></RESULT><RESULT eventid="32" heatid="346" lane="5" points="127" resultid="2579" swimtime="00:01:53.02"><SPLITS><SPLIT distance="50" swimtime="00:00:53.68"/></SPLITS></RESULT><RESULT eventid="36" heatid="384" lane="6" points="59" resultid="2860" swimtime="00:00:57.09"><SPLITS/></RESULT><RESULT eventid="38" heatid="414" lane="5" points="180" resultid="3087" swimtime="00:03:18.17"><SPLITS><SPLIT distance="50" swimtime="00:00:47.03"/><SPLIT distance="100" swimtime="00:01:37.40"/><SPLIT distance="150" swimtime="00:02:29.04"/></SPLITS></RESULT><RESULT eventid="40" heatid="453" lane="1" points="136" resultid="3382" swimtime="00:01:31.00"><SPLITS><SPLIT distance="50" swimtime="00:00:43.49"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="535" birthdate="2012-01-01" firstname="Myroslav" gender="M" lastname="Mymrenko" license="504586"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="10" heatid="132" lane="3" points="130" resultid="997" swimtime="00:00:41.24"><SPLITS/></RESULT><RESULT eventid="28" heatid="273" lane="7" points="137" resultid="2030" swimtime="00:00:45.92"><SPLITS/></RESULT><RESULT eventid="40" heatid="451" lane="5" points="102" resultid="3370" swimtime="00:01:40.28"><SPLITS><SPLIT distance="50" swimtime="00:00:43.17"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="537" birthdate="2010-01-01" firstname="Hannes" gender="M" lastname="Jannack" license="504315"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="10" heatid="132" lane="5" points="230" resultid="999" swimtime="00:00:34.12"><SPLITS/></RESULT><RESULT eventid="28" heatid="273" lane="2" points="185" resultid="2025" swimtime="00:00:41.57"><SPLITS/></RESULT><RESULT eventid="30" heatid="308" lane="4" points="202" resultid="2293" swimtime="00:02:53.71"><SPLITS><SPLIT distance="50" swimtime="00:00:37.30"/><SPLIT distance="100" swimtime="00:01:20.90"/><SPLIT distance="150" swimtime="00:02:06.52"/></SPLITS></RESULT><RESULT eventid="40" heatid="451" lane="8" points="220" resultid="3373" swimtime="00:01:17.60"><SPLITS><SPLIT distance="50" swimtime="00:00:37.21"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="538" birthdate="2012-01-01" firstname="Timofei" gender="M" lastname="Tsvetkov" license="504658"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="10" heatid="133" lane="7" points="95" resultid="1005" swimtime="00:00:45.80"><SPLITS/></RESULT><RESULT eventid="40" heatid="451" lane="6" points="87" resultid="3371" swimtime="00:01:45.54"><SPLITS><SPLIT distance="50" swimtime="00:00:46.94"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="539" birthdate="2016-01-01" firstname="Luka" gender="M" lastname="Lazic" license="499226"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="10" heatid="134" lane="2" points="105" resultid="1007" swimtime="00:00:44.30"><SPLITS/></RESULT><RESULT eventid="14" heatid="211" lane="8" points="99" resultid="1604" swimtime="00:01:51.21"><SPLITS><SPLIT distance="50" swimtime="00:00:53.74"/></SPLITS></RESULT><RESULT eventid="28" heatid="274" lane="3" points="85" resultid="2033" swimtime="00:00:53.90"><SPLITS/></RESULT><RESULT eventid="30" heatid="309" lane="2" points="82" resultid="2297" swimtime="00:03:54.00"><SPLITS><SPLIT distance="50" swimtime="00:00:53.99"/><SPLIT distance="100" swimtime="00:01:55.62"/><SPLIT distance="150" swimtime="00:02:58.83"/></SPLITS></RESULT><RESULT eventid="40" heatid="452" lane="4" points="80" resultid="3377" swimtime="00:01:48.34"><SPLITS><SPLIT distance="50" swimtime="00:00:53.56"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="540" birthdate="2016-01-01" firstname="Ilhan" gender="M" lastname="Yesilbag" license="498417"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="10" heatid="135" lane="8" points="73" resultid="1020" swimtime="00:00:49.85"><SPLITS/></RESULT><RESULT eventid="14" heatid="210" lane="5" points="108" resultid="1594" swimtime="00:01:48.03"><SPLITS><SPLIT distance="50" swimtime="00:00:52.25"/></SPLITS></RESULT><RESULT eventid="28" heatid="277" lane="8" points="100" resultid="2060" swimtime="00:00:50.98"><SPLITS/></RESULT><RESULT eventid="30" heatid="309" lane="3" points="82" resultid="2298" swimtime="00:03:54.72"><SPLITS><SPLIT distance="50" swimtime="00:00:53.93"/><SPLIT distance="100" swimtime="00:01:56.16"/><SPLIT distance="150" swimtime="00:02:59.55"/></SPLITS></RESULT><RESULT eventid="40" heatid="452" lane="6" points="67" resultid="3379" swimtime="00:01:55.01"><SPLITS><SPLIT distance="50" swimtime="00:00:54.59"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="572" birthdate="2016-01-01" firstname="Aurora" gender="F" lastname="Busse" license="495895"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="27" heatid="254" lane="7" points="78" resultid="1882" swimtime="00:01:03.07"><SPLITS/></RESULT><RESULT eventid="31" heatid="328" lane="4" points="152" resultid="2438" swimtime="00:02:00.09"><SPLITS><SPLIT distance="50" swimtime="00:00:57.86"/></SPLITS></RESULT><RESULT eventid="39" heatid="420" lane="4" points="78" resultid="3128" swimtime="00:02:00.82"><SPLITS><SPLIT distance="50" swimtime="00:00:54.82"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="588" birthdate="2016-01-01" firstname="Abaan" gender="M" lastname="Khan" license="504320"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="28" heatid="273" lane="4" points="27" resultid="2027" swimtime="00:01:18.30"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="589" birthdate="2011-01-01" firstname="Niklas" gender="M" lastname="Blumhagen" license="504306"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="28" heatid="273" lane="5" points="115" resultid="2028" swimtime="00:00:48.62"><SPLITS/></RESULT><RESULT eventid="30" heatid="308" lane="3" points="98" resultid="2292" swimtime="00:03:40.66"><SPLITS><SPLIT distance="50" swimtime="00:00:45.24"/><SPLIT distance="100" swimtime="00:01:43.38"/><SPLIT distance="150" swimtime="00:02:44.02"/></SPLITS></RESULT><RESULT eventid="32" heatid="345" lane="4" points="147" resultid="2572" swimtime="00:01:47.65"><SPLITS><SPLIT distance="50" swimtime="00:00:48.54"/></SPLITS></RESULT><RESULT eventid="40" heatid="452" lane="8" points="110" resultid="3381" swimtime="00:01:37.51"><SPLITS><SPLIT distance="50" swimtime="00:00:45.01"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="590" birthdate="2013-01-01" firstname="Manuel" gender="M" lastname="Blumhagen" license="504305"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="28" heatid="273" lane="6" points="52" resultid="2029" swimtime="00:01:03.38"><SPLITS/></RESULT><RESULT eventid="32" heatid="345" lane="5" points="97" resultid="2573" swimtime="00:02:03.74"><SPLITS><SPLIT distance="50" swimtime="00:00:57.56"/></SPLITS></RESULT><RESULT eventid="40" heatid="451" lane="4" points="44" resultid="3369" swimtime="00:02:12.49"><SPLITS><SPLIT distance="50" swimtime="00:00:58.57"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="605" birthdate="2012-01-01" firstname="Roman" gender="M" lastname="Shevchenko" license="504317"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="32" heatid="345" lane="6" points="128" resultid="2574" swimtime="00:01:52.78"><SPLITS><SPLIT distance="50" swimtime="00:00:52.24"/></SPLITS></RESULT><RESULT eventid="40" heatid="451" lane="1" points="124" resultid="3366" swimtime="00:01:33.75"><SPLITS><SPLIT distance="50" swimtime="00:00:40.92"/></SPLITS></RESULT></RESULTS></ATHLETE></ATHLETES><RELAYS/></CLUB><CLUB code="4958" name="SSG 81 Erlangen" nation="GER" region="02" shortname="Erlangen" type="CLUB"><CONTACT city="Erlangen" country="GER" email="roland.boeller@gmx.de" name="Böller, Roland" phone="0178/1606404" street="Adalbert-Stifter-Str. 8" zip="91054"/><OFFICIALS/><ATHLETES><ATHLETE athleteid="9" birthdate="2016-01-01" firstname="Dana" gender="F" lastname="Puchalla" license="491822"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="2" lane="5" points="72" resultid="9" swimtime="00:01:10.14"><SPLITS/></RESULT><RESULT eventid="9" heatid="103" lane="5" points="100" resultid="773" swimtime="00:00:50.85"><SPLITS/></RESULT><RESULT eventid="27" heatid="253" lane="2" points="94" resultid="1869" swimtime="00:00:59.17"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="13" birthdate="2016-01-01" firstname="Lara" gender="F" lastname="Schenk" license="491157"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="3" lane="1" points="85" resultid="13" swimtime="00:01:06.52"><SPLITS/></RESULT><RESULT eventid="9" heatid="104" lane="8" points="87" resultid="784" swimtime="00:00:53.31"><SPLITS/></RESULT><RESULT eventid="27" heatid="254" lane="3" points="114" resultid="1878" swimtime="00:00:55.61"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="15" birthdate="2013-01-01" firstname="Julia" gender="F" lastname="Kurth" license="462967"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="3" lane="3" points="117" resultid="15" swimtime="00:00:59.87"><SPLITS/></RESULT><RESULT eventid="9" heatid="106" lane="5" points="131" resultid="797" swimtime="00:00:46.60"><SPLITS/></RESULT><RESULT eventid="13" heatid="191" lane="6" points="138" resultid="1445" swimtime="00:01:50.94"><SPLITS><SPLIT distance="50" swimtime="00:00:51.43"/></SPLITS></RESULT><RESULT eventid="27" heatid="257" lane="2" points="149" resultid="1901" swimtime="00:00:50.87"><SPLITS/></RESULT><RESULT eventid="31" heatid="327" lane="5" points="116" resultid="2432" swimtime="00:02:11.27"><SPLITS><SPLIT distance="50" swimtime="00:01:00.92"/></SPLITS></RESULT><RESULT eventid="35" heatid="363" lane="2" points="61" resultid="2697" swimtime="00:01:01.73"><SPLITS/></RESULT><RESULT eventid="39" heatid="422" lane="4" points="120" resultid="3142" swimtime="00:01:44.67"><SPLITS><SPLIT distance="50" swimtime="00:00:49.64"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="27" birthdate="2014-01-01" firstname="Ronja" gender="F" lastname="Kurth" license="462968"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="4" lane="7" points="149" resultid="27" swimtime="00:00:55.18"><SPLITS/></RESULT><RESULT eventid="9" heatid="111" lane="6" points="222" resultid="838" swimtime="00:00:39.08"><SPLITS/></RESULT><RESULT eventid="13" heatid="192" lane="8" points="136" resultid="1455" swimtime="00:01:51.57"><SPLITS><SPLIT distance="50" swimtime="00:00:54.15"/></SPLITS></RESULT><RESULT eventid="27" heatid="257" lane="6" points="151" resultid="1905" swimtime="00:00:50.56"><SPLITS/></RESULT><RESULT eventid="29" heatid="290" lane="8" points="148" resultid="2158" swimtime="00:03:33.31"><SPLITS><SPLIT distance="50" swimtime="00:00:47.91"/><SPLIT distance="100" swimtime="00:01:43.19"/><SPLIT distance="150" swimtime="00:02:40.97"/></SPLITS></RESULT><RESULT eventid="31" heatid="328" lane="8" points="159" resultid="2442" swimtime="00:01:58.26"><SPLITS><SPLIT distance="50" swimtime="00:00:59.05"/></SPLITS></RESULT><RESULT eventid="35" heatid="363" lane="5" points="78" resultid="2699" swimtime="00:00:57.00"><SPLITS/></RESULT><RESULT eventid="39" heatid="426" lane="8" resultid="3177" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="30" birthdate="2015-01-01" firstname="Joana" gender="F" lastname="Kojro" license="479247"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="5" lane="2" points="148" resultid="30" swimtime="00:00:55.34"><SPLITS/></RESULT><RESULT eventid="3" heatid="46" lane="8" points="329" resultid="351" swimtime="00:05:42.38"><SPLITS><SPLIT distance="100" swimtime="00:01:20.91"/><SPLIT distance="200" swimtime="00:02:49.13"/><SPLIT distance="300" swimtime="00:04:18.73"/></SPLITS></RESULT><RESULT eventid="9" heatid="114" lane="4" points="305" resultid="860" swimtime="00:00:35.16"><SPLITS/></RESULT><RESULT eventid="11" heatid="160" lane="7" points="238" resultid="1209" swimtime="00:03:23.37"><SPLITS><SPLIT distance="50" swimtime="00:00:48.18"/><SPLIT distance="100" swimtime="00:01:35.60"/><SPLIT distance="150" swimtime="00:02:41.56"/></SPLITS></RESULT><RESULT eventid="27" heatid="262" lane="8" points="252" resultid="1947" swimtime="00:00:42.66"><SPLITS/></RESULT><RESULT eventid="29" heatid="296" lane="6" points="348" resultid="2203" swimtime="00:02:40.51"><SPLITS><SPLIT distance="50" swimtime="00:00:37.36"/><SPLIT distance="100" swimtime="00:01:19.25"/><SPLIT distance="150" swimtime="00:02:00.34"/></SPLITS></RESULT><RESULT eventid="35" heatid="368" lane="3" points="175" resultid="2737" swimtime="00:00:43.63"><SPLITS/></RESULT><RESULT eventid="39" heatid="434" lane="1" points="304" resultid="3234" swimtime="00:01:16.86"><SPLITS><SPLIT distance="50" swimtime="00:00:37.52"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="44" birthdate="2014-01-01" firstname="Lisa" gender="F" lastname="Hahn" license="479759"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="6" lane="8" points="126" resultid="44" swimtime="00:00:58.33"><SPLITS/></RESULT><RESULT eventid="9" heatid="108" lane="3" points="154" resultid="811" swimtime="00:00:44.14"><SPLITS/></RESULT><RESULT eventid="13" heatid="190" lane="2" points="91" resultid="1435" swimtime="00:02:07.54"><SPLITS><SPLIT distance="50" swimtime="00:00:59.77"/></SPLITS></RESULT><RESULT eventid="27" heatid="255" lane="7" points="133" resultid="1890" swimtime="00:00:52.74"><SPLITS/></RESULT><RESULT eventid="31" heatid="328" lane="1" points="143" resultid="2435" swimtime="00:02:02.37"><SPLITS><SPLIT distance="50" swimtime="00:01:01.10"/></SPLITS></RESULT><RESULT eventid="39" heatid="421" lane="2" points="125" resultid="3132" swimtime="00:01:43.22"><SPLITS><SPLIT distance="50" swimtime="00:00:49.47"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="46" birthdate="2014-01-01" firstname="Ezgi" gender="F" lastname="Özden" license="462888"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="7" lane="2" points="163" resultid="46" swimtime="00:00:53.54"><SPLITS/></RESULT><RESULT eventid="9" heatid="107" lane="4" points="183" resultid="804" swimtime="00:00:41.62"><SPLITS/></RESULT><RESULT eventid="13" heatid="194" lane="2" points="144" resultid="1465" swimtime="00:01:49.38"><SPLITS><SPLIT distance="50" swimtime="00:00:51.08"/></SPLITS></RESULT><RESULT eventid="27" heatid="258" lane="1" points="167" resultid="1908" swimtime="00:00:48.92"><SPLITS/></RESULT><RESULT eventid="31" heatid="328" lane="7" points="175" resultid="2441" swimtime="00:01:54.65"><SPLITS><SPLIT distance="50" swimtime="00:00:54.54"/></SPLITS></RESULT><RESULT eventid="35" heatid="364" lane="3" points="111" resultid="2705" swimtime="00:00:50.83"><SPLITS/></RESULT><RESULT eventid="39" heatid="423" lane="1" points="139" resultid="3147" swimtime="00:01:39.65"><SPLITS><SPLIT distance="50" swimtime="00:00:49.26"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="50" birthdate="2015-01-01" firstname="Cara Luna" gender="F" lastname="Burnes" license="476018"><HANDICAP/><ENTRIES/><RESULTS><RESULT comment="09:18 Start vor dem Startsignal" eventid="1" heatid="7" lane="6" resultid="50" status="DSQ" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="9" heatid="105" lane="1" points="145" resultid="785" swimtime="00:00:44.98"><SPLITS/></RESULT><RESULT eventid="13" heatid="191" lane="2" points="126" resultid="1441" swimtime="00:01:54.52"><SPLITS><SPLIT distance="50" swimtime="00:00:51.91"/></SPLITS></RESULT><RESULT eventid="27" heatid="254" lane="4" points="130" resultid="1879" swimtime="00:00:53.20"><SPLITS/></RESULT><RESULT eventid="39" heatid="421" lane="6" points="114" resultid="3136" swimtime="00:01:46.62"><SPLITS><SPLIT distance="50" swimtime="00:00:48.64"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="58" birthdate="2013-01-01" firstname="Malak" gender="F" lastname="Khalil" license="489783"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="8" lane="6" points="185" resultid="58" swimtime="00:00:51.40"><SPLITS/></RESULT><RESULT eventid="9" heatid="108" lane="5" points="160" resultid="813" swimtime="00:00:43.52"><SPLITS/></RESULT><RESULT eventid="25" heatid="247" lane="7" resultid="1836" swimtime="00:01:00.90"><SPLITS/></RESULT><RESULT eventid="31" heatid="331" lane="8" points="175" resultid="2466" swimtime="00:01:54.45"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="67" birthdate="2014-01-01" firstname="Josephine Alexia" gender="F" lastname="Baker-Duly" license="460130"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="9" lane="7" points="163" resultid="67" swimtime="00:00:53.60"><SPLITS/></RESULT><RESULT eventid="9" heatid="110" lane="4" points="221" resultid="828" swimtime="00:00:39.14"><SPLITS/></RESULT><RESULT eventid="13" heatid="193" lane="2" points="160" resultid="1457" swimtime="00:01:45.66"><SPLITS><SPLIT distance="50" swimtime="00:00:52.83"/></SPLITS></RESULT><RESULT eventid="27" heatid="257" lane="8" points="138" resultid="1907" swimtime="00:00:52.18"><SPLITS/></RESULT><RESULT eventid="31" heatid="331" lane="6" points="182" resultid="2464" swimtime="00:01:53.03"><SPLITS/></RESULT><RESULT eventid="39" heatid="427" lane="4" points="188" resultid="3181" swimtime="00:01:30.25"><SPLITS><SPLIT distance="50" swimtime="00:00:44.16"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="70" birthdate="2013-01-01" firstname="Wanying" gender="F" lastname="Sun" license="470922"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="10" lane="2" points="174" resultid="70" swimtime="00:00:52.47"><SPLITS/></RESULT><RESULT eventid="7" heatid="83" lane="1" points="187" resultid="618" swimtime="00:04:02.78"><SPLITS><SPLIT distance="50" swimtime="00:00:54.97"/><SPLIT distance="100" swimtime="00:01:57.43"/><SPLIT distance="150" swimtime="00:03:01.30"/></SPLITS></RESULT><RESULT eventid="9" heatid="111" lane="2" points="221" resultid="834" swimtime="00:00:39.13"><SPLITS/></RESULT><RESULT eventid="11" heatid="159" lane="8" points="168" resultid="1202" swimtime="00:03:48.13"><SPLITS><SPLIT distance="50" swimtime="00:00:55.85"/><SPLIT distance="100" swimtime="00:01:51.70"/><SPLIT distance="150" swimtime="00:02:57.83"/></SPLITS></RESULT><RESULT eventid="29" heatid="292" lane="5" points="212" resultid="2170" swimtime="00:03:09.21"><SPLITS><SPLIT distance="50" swimtime="00:00:44.01"/><SPLIT distance="100" swimtime="00:01:32.68"/><SPLIT distance="150" swimtime="00:02:23.21"/></SPLITS></RESULT><RESULT eventid="31" heatid="332" lane="6" points="175" resultid="2472" swimtime="00:01:54.47"><SPLITS><SPLIT distance="50" swimtime="00:00:54.77"/></SPLITS></RESULT><RESULT eventid="39" heatid="429" lane="3" points="204" resultid="3196" swimtime="00:01:27.72"><SPLITS><SPLIT distance="50" swimtime="00:00:43.89"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="71" birthdate="2015-01-01" firstname="Céline" gender="F" lastname="Ettinger" license="460135"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="10" lane="3" points="176" resultid="71" swimtime="00:00:52.20"><SPLITS/></RESULT><RESULT eventid="9" heatid="111" lane="3" points="253" resultid="835" swimtime="00:00:37.39"><SPLITS/></RESULT><RESULT eventid="13" heatid="196" lane="6" points="177" resultid="1485" swimtime="00:01:42.21"><SPLITS><SPLIT distance="50" swimtime="00:00:45.84"/></SPLITS></RESULT><RESULT eventid="27" heatid="260" lane="8" resultid="1931" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="31" heatid="331" lane="1" resultid="2459" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="39" heatid="427" lane="5" resultid="3182" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="75" birthdate="2013-01-01" firstname="Hannah" gender="F" lastname="Lechler" license="478966"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="10" lane="7" points="165" resultid="75" swimtime="00:00:53.34"><SPLITS/></RESULT><RESULT eventid="9" heatid="109" lane="3" points="172" resultid="819" swimtime="00:00:42.48"><SPLITS/></RESULT><RESULT eventid="27" heatid="256" lane="3" points="155" resultid="1894" swimtime="00:00:50.22"><SPLITS/></RESULT><RESULT eventid="29" heatid="289" lane="1" points="103" resultid="2143" swimtime="00:04:00.73"><SPLITS><SPLIT distance="50" swimtime="00:00:47.89"/><SPLIT distance="100" swimtime="00:01:47.84"/><SPLIT distance="150" swimtime="00:02:56.21"/></SPLITS></RESULT><RESULT eventid="31" heatid="329" lane="8" points="156" resultid="2450" swimtime="00:01:59.01"><SPLITS><SPLIT distance="50" swimtime="00:00:56.63"/></SPLITS></RESULT><RESULT eventid="35" heatid="363" lane="6" points="66" resultid="2700" swimtime="00:01:00.26"><SPLITS/></RESULT><RESULT eventid="39" heatid="424" lane="4" points="137" resultid="3158" swimtime="00:01:40.14"><SPLITS><SPLIT distance="50" swimtime="00:00:47.38"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="76" birthdate="2014-01-01" firstname="Lisa" gender="F" lastname="Schenk" license="460205"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="10" lane="8" points="171" resultid="76" swimtime="00:00:52.69"><SPLITS/></RESULT><RESULT eventid="7" heatid="83" lane="2" points="210" resultid="619" swimtime="00:03:53.42"><SPLITS><SPLIT distance="50" swimtime="00:00:54.51"/><SPLIT distance="100" swimtime="00:01:51.84"/><SPLIT distance="150" swimtime="00:02:53.65"/></SPLITS></RESULT><RESULT eventid="9" heatid="107" lane="8" points="130" resultid="808" swimtime="00:00:46.69"><SPLITS/></RESULT><RESULT eventid="27" heatid="255" lane="4" points="104" resultid="1887" swimtime="00:00:57.28"><SPLITS/></RESULT><RESULT eventid="31" heatid="332" lane="4" points="187" resultid="2470" swimtime="00:01:51.97"><SPLITS><SPLIT distance="50" swimtime="00:00:52.96"/></SPLITS></RESULT><RESULT eventid="39" heatid="424" lane="8" points="115" resultid="3162" swimtime="00:01:46.10"><SPLITS><SPLIT distance="50" swimtime="00:00:49.87"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="79" birthdate="2014-01-01" firstname="Sofiia" gender="F" lastname="Lukina" license="470855"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="11" lane="3" points="223" resultid="79" swimtime="00:00:48.31"><SPLITS/></RESULT><RESULT eventid="7" heatid="84" lane="3" points="239" resultid="627" swimtime="00:03:43.64"><SPLITS><SPLIT distance="50" swimtime="00:00:51.48"/><SPLIT distance="100" swimtime="00:01:49.49"/><SPLIT distance="150" swimtime="00:02:47.56"/></SPLITS></RESULT><RESULT eventid="9" heatid="113" lane="8" points="226" resultid="856" swimtime="00:00:38.83"><SPLITS/></RESULT><RESULT eventid="13" heatid="195" lane="4" points="206" resultid="1475" swimtime="00:01:37.27"><SPLITS><SPLIT distance="50" swimtime="00:00:47.35"/></SPLITS></RESULT><RESULT eventid="27" heatid="259" lane="2" points="218" resultid="1917" swimtime="00:00:44.80"><SPLITS/></RESULT><RESULT eventid="29" heatid="293" lane="2" points="250" resultid="2175" swimtime="00:02:59.29"><SPLITS><SPLIT distance="50" swimtime="00:00:42.39"/><SPLIT distance="100" swimtime="00:01:28.44"/><SPLIT distance="150" swimtime="00:02:15.68"/></SPLITS></RESULT><RESULT eventid="35" heatid="366" lane="1" points="128" resultid="2719" swimtime="00:00:48.43"><SPLITS/></RESULT><RESULT eventid="39" heatid="428" lane="6" points="240" resultid="3191" swimtime="00:01:23.10"><SPLITS><SPLIT distance="50" swimtime="00:00:41.21"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="85" birthdate="2012-01-01" firstname="Iuliia" gender="F" lastname="Kazakova" license="479355"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="12" lane="1" points="218" resultid="85" swimtime="00:00:48.67"><SPLITS/></RESULT><RESULT eventid="9" heatid="119" lane="8" points="383" resultid="903" swimtime="00:00:32.58"><SPLITS/></RESULT><RESULT eventid="13" heatid="196" lane="2" points="317" resultid="1481" swimtime="00:01:24.22"><SPLITS><SPLIT distance="50" swimtime="00:00:42.03"/></SPLITS></RESULT><RESULT eventid="27" heatid="263" lane="3" points="335" resultid="1950" swimtime="00:00:38.82"><SPLITS/></RESULT><RESULT eventid="29" heatid="300" lane="8" points="354" resultid="2237" swimtime="00:02:39.59"><SPLITS><SPLIT distance="50" swimtime="00:00:36.81"/><SPLIT distance="100" swimtime="00:01:17.24"/><SPLIT distance="150" swimtime="00:02:00.31"/></SPLITS></RESULT><RESULT eventid="35" heatid="372" lane="1" points="263" resultid="2767" swimtime="00:00:38.11"><SPLITS/></RESULT><RESULT eventid="39" heatid="436" lane="4" points="344" resultid="3253" swimtime="00:01:13.77"><SPLITS><SPLIT distance="50" swimtime="00:00:35.81"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="90" birthdate="2013-01-01" firstname="Frida Adelaide" gender="F" lastname="Baker-Duly" license="460129"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="12" lane="6" points="260" resultid="90" swimtime="00:00:45.86"><SPLITS/></RESULT><RESULT eventid="7" heatid="85" lane="6" points="261" resultid="638" swimtime="00:03:37.17"><SPLITS><SPLIT distance="50" swimtime="00:00:49.09"/><SPLIT distance="100" swimtime="00:01:44.78"/><SPLIT distance="150" swimtime="00:02:41.85"/></SPLITS></RESULT><RESULT eventid="9" heatid="112" lane="8" points="209" resultid="848" swimtime="00:00:39.84"><SPLITS/></RESULT><RESULT eventid="31" heatid="337" lane="1" points="248" resultid="2507" swimtime="00:01:42.02"><SPLITS><SPLIT distance="50" swimtime="00:00:49.24"/></SPLITS></RESULT><RESULT eventid="35" heatid="366" lane="8" points="117" resultid="2726" swimtime="00:00:49.89"><SPLITS/></RESULT><RESULT eventid="39" heatid="429" lane="5" points="191" resultid="3198" swimtime="00:01:29.76"><SPLITS><SPLIT distance="50" swimtime="00:00:44.05"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="93" birthdate="2009-01-01" firstname="Viktoria" gender="F" lastname="Biró" license="409145"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="13" lane="1" points="199" resultid="93" swimtime="00:00:50.17"><SPLITS/></RESULT><RESULT eventid="9" heatid="116" lane="5" points="289" resultid="877" swimtime="00:00:35.79"><SPLITS/></RESULT><RESULT eventid="13" heatid="200" lane="3" points="310" resultid="1514" swimtime="00:01:24.84"><SPLITS/></RESULT><RESULT eventid="29" heatid="296" lane="4" points="296" resultid="2201" swimtime="00:02:49.51"><SPLITS><SPLIT distance="50" swimtime="00:00:37.95"/><SPLIT distance="100" swimtime="00:01:21.00"/><SPLIT distance="150" swimtime="00:02:06.18"/></SPLITS></RESULT><RESULT eventid="35" heatid="369" lane="1" points="156" resultid="2743" swimtime="00:00:45.31"><SPLITS/></RESULT><RESULT eventid="39" heatid="434" lane="8" points="260" resultid="3241" swimtime="00:01:20.96"><SPLITS><SPLIT distance="50" swimtime="00:00:39.81"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="94" birthdate="2009-01-01" firstname="Anna Helene" gender="F" lastname="Richter" license="409131"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="13" lane="2" points="241" resultid="94" swimtime="00:00:47.04"><SPLITS/></RESULT><RESULT eventid="9" heatid="114" lane="6" points="273" resultid="862" swimtime="00:00:36.45"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="95" birthdate="2016-01-01" firstname="Marie" gender="F" lastname="Marschall" license="479176"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="13" lane="3" points="214" resultid="95" swimtime="00:00:48.97"><SPLITS/></RESULT><RESULT eventid="9" heatid="114" lane="1" points="228" resultid="857" swimtime="00:00:38.72"><SPLITS/></RESULT><RESULT eventid="27" heatid="259" lane="1" points="204" resultid="1916" swimtime="00:00:45.79"><SPLITS/></RESULT><RESULT eventid="29" heatid="293" lane="6" points="202" resultid="2179" swimtime="00:03:12.48"><SPLITS><SPLIT distance="50" swimtime="00:00:41.09"/><SPLIT distance="100" swimtime="00:01:31.16"/><SPLIT distance="150" swimtime="00:02:23.45"/></SPLITS></RESULT><RESULT eventid="35" heatid="365" lane="4" points="133" resultid="2714" swimtime="00:00:47.80"><SPLITS/></RESULT><RESULT eventid="39" heatid="430" lane="1" points="231" resultid="3202" swimtime="00:01:24.22"><SPLITS><SPLIT distance="50" swimtime="00:00:39.61"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="98" birthdate="2013-01-01" firstname="Julia" gender="F" lastname="Neugebauer" license="460203"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="13" lane="6" points="224" resultid="98" swimtime="00:00:48.22"><SPLITS/></RESULT><RESULT eventid="9" heatid="114" lane="5" points="290" resultid="861" swimtime="00:00:35.74"><SPLITS/></RESULT><RESULT eventid="13" heatid="198" lane="6" points="192" resultid="1501" swimtime="00:01:39.42"><SPLITS><SPLIT distance="50" swimtime="00:00:50.04"/></SPLITS></RESULT><RESULT eventid="27" heatid="261" lane="2" points="216" resultid="1933" swimtime="00:00:44.96"><SPLITS/></RESULT><RESULT eventid="31" heatid="335" lane="6" points="231" resultid="2496" swimtime="00:01:44.41"><SPLITS><SPLIT distance="50" swimtime="00:00:50.32"/></SPLITS></RESULT><RESULT eventid="39" heatid="430" lane="7" points="226" resultid="3208" swimtime="00:01:24.88"><SPLITS><SPLIT distance="50" swimtime="00:00:41.51"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="100" birthdate="2011-01-01" firstname="Sophie" gender="F" lastname="Henglein" license="447064"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="13" lane="8" points="216" resultid="100" swimtime="00:00:48.78"><SPLITS/></RESULT><RESULT eventid="9" heatid="112" lane="2" points="319" resultid="842" swimtime="00:00:34.64"><SPLITS/></RESULT><RESULT eventid="11" heatid="159" lane="1" points="240" resultid="1196" swimtime="00:03:22.72"><SPLITS><SPLIT distance="50" swimtime="00:00:46.58"/><SPLIT distance="100" swimtime="00:01:37.55"/><SPLIT distance="150" swimtime="00:02:38.25"/></SPLITS></RESULT><RESULT eventid="27" heatid="256" lane="4" points="213" resultid="1895" swimtime="00:00:45.16"><SPLITS/></RESULT><RESULT eventid="31" heatid="335" lane="5" points="215" resultid="2495" swimtime="00:01:47.00"><SPLITS><SPLIT distance="50" swimtime="00:00:50.13"/></SPLITS></RESULT><RESULT eventid="35" heatid="367" lane="2" points="201" resultid="2728" swimtime="00:00:41.66"><SPLITS/></RESULT><RESULT eventid="39" heatid="431" lane="4" points="273" resultid="3213" swimtime="00:01:19.68"><SPLITS><SPLIT distance="50" swimtime="00:00:36.73"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="101" birthdate="2013-01-01" firstname="Emilia" gender="F" lastname="Häring" license="462955"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="14" lane="1" resultid="101" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="27" heatid="258" lane="7" resultid="1914" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="29" heatid="289" lane="3" resultid="2145" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="31" heatid="334" lane="6" resultid="2488" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="39" heatid="426" lane="4" resultid="3173" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="104" birthdate="2011-01-01" firstname="Carolina" gender="F" lastname="Beyfuß" license="446470"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="14" lane="4" points="255" resultid="104" swimtime="00:00:46.20"><SPLITS/></RESULT><RESULT eventid="7" heatid="86" lane="7" points="259" resultid="647" swimtime="00:03:37.87"><SPLITS><SPLIT distance="50" swimtime="00:00:49.22"/><SPLIT distance="100" swimtime="00:01:44.87"/><SPLIT distance="150" swimtime="00:02:43.71"/></SPLITS></RESULT><RESULT eventid="9" heatid="112" lane="5" points="260" resultid="845" swimtime="00:00:37.07"><SPLITS/></RESULT><RESULT eventid="13" heatid="196" lane="4" points="230" resultid="1483" swimtime="00:01:33.70"><SPLITS><SPLIT distance="50" swimtime="00:00:44.21"/></SPLITS></RESULT><RESULT eventid="29" heatid="295" lane="3" points="244" resultid="2192" swimtime="00:03:00.59"><SPLITS><SPLIT distance="50" swimtime="00:00:40.45"/><SPLIT distance="100" swimtime="00:01:26.03"/><SPLIT distance="150" swimtime="00:02:14.98"/></SPLITS></RESULT><RESULT eventid="35" heatid="367" lane="5" points="197" resultid="2731" swimtime="00:00:41.97"><SPLITS/></RESULT><RESULT eventid="39" heatid="432" lane="1" points="251" resultid="3218" swimtime="00:01:21.90"><SPLITS><SPLIT distance="50" swimtime="00:00:39.91"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="108" birthdate="2015-01-01" firstname="Leni" gender="F" lastname="Moosmeier" license="470675"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="14" lane="8" points="244" resultid="108" swimtime="00:00:46.83"><SPLITS/></RESULT><RESULT eventid="7" heatid="86" lane="2" points="264" resultid="642" swimtime="00:03:36.40"><SPLITS><SPLIT distance="50" swimtime="00:00:50.09"/><SPLIT distance="100" swimtime="00:01:45.41"/><SPLIT distance="150" swimtime="00:02:43.45"/></SPLITS></RESULT><RESULT eventid="11" heatid="161" lane="5" points="254" resultid="1215" swimtime="00:03:19.01"><SPLITS><SPLIT distance="50" swimtime="00:00:44.07"/><SPLIT distance="100" swimtime="00:01:39.94"/><SPLIT distance="150" swimtime="00:02:36.52"/></SPLITS></RESULT><RESULT eventid="13" heatid="199" lane="2" points="192" resultid="1505" swimtime="00:01:39.45"><SPLITS><SPLIT distance="50" swimtime="00:00:48.99"/></SPLITS></RESULT><RESULT eventid="29" heatid="290" lane="4" points="266" resultid="2154" swimtime="00:02:55.67"><SPLITS><SPLIT distance="50" swimtime="00:00:39.43"/><SPLIT distance="100" swimtime="00:01:24.72"/><SPLIT distance="150" swimtime="00:02:11.17"/></SPLITS></RESULT><RESULT eventid="31" heatid="335" lane="4" points="236" resultid="2494" swimtime="00:01:43.74"><SPLITS><SPLIT distance="50" swimtime="00:00:49.79"/></SPLITS></RESULT><RESULT eventid="35" heatid="368" lane="4" points="178" resultid="2738" swimtime="00:00:43.36"><SPLITS/></RESULT><RESULT eventid="39" heatid="426" lane="6" points="257" resultid="3175" swimtime="00:01:21.27"><SPLITS><SPLIT distance="50" swimtime="00:00:38.51"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="115" birthdate="2013-01-01" firstname="Carlotta" gender="F" lastname="Stein" license="450788"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="15" lane="7" points="224" resultid="115" swimtime="00:00:48.24"><SPLITS/></RESULT><RESULT eventid="5" heatid="65" lane="6" points="276" resultid="486" swimtime="00:01:25.15"><SPLITS><SPLIT distance="50" swimtime="00:00:37.30"/></SPLITS></RESULT><RESULT eventid="9" heatid="117" lane="3" points="310" resultid="882" swimtime="00:00:34.95"><SPLITS/></RESULT><RESULT eventid="11" heatid="165" lane="1" points="303" resultid="1243" swimtime="00:03:07.72"><SPLITS><SPLIT distance="50" swimtime="00:00:41.28"/><SPLIT distance="100" swimtime="00:01:30.72"/><SPLIT distance="150" swimtime="00:02:25.62"/></SPLITS></RESULT><RESULT eventid="27" heatid="267" lane="3" points="340" resultid="1982" swimtime="00:00:38.63"><SPLITS/></RESULT><RESULT eventid="31" heatid="330" lane="3" points="229" resultid="2453" swimtime="00:01:44.73"><SPLITS/></RESULT><RESULT eventid="35" heatid="372" lane="5" points="282" resultid="2771" swimtime="00:00:37.24"><SPLITS/></RESULT><RESULT eventid="39" heatid="435" lane="4" points="295" resultid="3245" swimtime="00:01:17.61"><SPLITS><SPLIT distance="50" swimtime="00:00:36.39"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="120" birthdate="2014-01-01" firstname="Nika" gender="F" lastname="Splihal" license="470857"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="16" lane="4" points="332" resultid="120" swimtime="00:00:42.31"><SPLITS/></RESULT><RESULT eventid="3" heatid="45" lane="3" points="280" resultid="338" swimtime="00:06:01.11"><SPLITS><SPLIT distance="100" swimtime="00:01:22.79"/><SPLIT distance="200" swimtime="00:02:55.72"/><SPLIT distance="300" swimtime="00:04:30.00"/></SPLITS></RESULT><RESULT eventid="7" heatid="87" lane="4" points="302" resultid="652" swimtime="00:03:27.03"><SPLITS><SPLIT distance="50" swimtime="00:00:45.96"/><SPLIT distance="100" swimtime="00:01:38.98"/><SPLIT distance="150" swimtime="00:02:34.04"/></SPLITS></RESULT><RESULT eventid="9" heatid="116" lane="7" points="300" resultid="879" swimtime="00:00:35.35"><SPLITS/></RESULT><RESULT eventid="11" heatid="163" lane="7" points="286" resultid="1233" swimtime="00:03:11.40"><SPLITS><SPLIT distance="50" swimtime="00:00:44.93"/><SPLIT distance="100" swimtime="00:01:34.10"/><SPLIT distance="150" swimtime="00:02:29.01"/></SPLITS></RESULT><RESULT eventid="25" heatid="249" lane="4" resultid="1848" swimtime="00:00:54.12"><SPLITS/></RESULT><RESULT eventid="31" heatid="337" lane="6" points="309" resultid="2512" swimtime="00:01:34.76"><SPLITS><SPLIT distance="50" swimtime="00:00:44.47"/></SPLITS></RESULT><RESULT eventid="39" heatid="435" lane="8" points="291" resultid="3249" swimtime="00:01:18.01"><SPLITS><SPLIT distance="50" swimtime="00:00:37.80"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="123" birthdate="2011-01-01" firstname="Ece" gender="F" lastname="Özden" license="446971"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="16" lane="7" points="247" resultid="123" swimtime="00:00:46.67"><SPLITS/></RESULT><RESULT eventid="5" heatid="63" lane="4" points="157" resultid="470" swimtime="00:01:42.63"><SPLITS><SPLIT distance="50" swimtime="00:00:46.11"/></SPLITS></RESULT><RESULT eventid="9" heatid="112" lane="6" points="259" resultid="846" swimtime="00:00:37.11"><SPLITS/></RESULT><RESULT eventid="27" heatid="259" lane="5" points="233" resultid="1920" swimtime="00:00:43.79"><SPLITS/></RESULT><RESULT eventid="31" heatid="336" lane="3" points="231" resultid="2501" swimtime="00:01:44.51"><SPLITS><SPLIT distance="50" swimtime="00:00:49.64"/></SPLITS></RESULT><RESULT eventid="35" heatid="367" lane="1" points="138" resultid="2727" swimtime="00:00:47.20"><SPLITS/></RESULT><RESULT eventid="39" heatid="430" lane="5" points="246" resultid="3206" swimtime="00:01:22.47"><SPLITS><SPLIT distance="50" swimtime="00:00:40.21"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="133" birthdate="2009-01-01" firstname="Hana" gender="F" lastname="Yaser Salih" license="404987"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="18" lane="1" resultid="133" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="9" heatid="116" lane="3" resultid="875" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="27" heatid="261" lane="1" resultid="1932" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="29" heatid="295" lane="8" resultid="2197" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="31" heatid="338" lane="5" resultid="2519" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="35" heatid="369" lane="8" resultid="2750" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="39" heatid="433" lane="2" resultid="3227" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="134" birthdate="2010-01-01" firstname="Dagrun" gender="F" lastname="Kraml" license="420928"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="18" lane="2" points="256" resultid="134" swimtime="00:00:46.12"><SPLITS/></RESULT><RESULT eventid="5" heatid="66" lane="5" points="250" resultid="493" swimtime="00:01:27.99"><SPLITS><SPLIT distance="50" swimtime="00:00:40.55"/></SPLITS></RESULT><RESULT eventid="9" heatid="120" lane="2" points="356" resultid="905" swimtime="00:00:33.39"><SPLITS/></RESULT><RESULT eventid="11" heatid="167" lane="2" points="282" resultid="1260" swimtime="00:03:12.25"><SPLITS><SPLIT distance="50" swimtime="00:00:38.66"/><SPLIT distance="100" swimtime="00:01:27.65"/><SPLIT distance="150" swimtime="00:02:23.29"/></SPLITS></RESULT><RESULT eventid="27" heatid="263" lane="7" points="287" resultid="1954" swimtime="00:00:40.86"><SPLITS/></RESULT><RESULT eventid="35" heatid="374" lane="5" points="284" resultid="2787" swimtime="00:00:37.15"><SPLITS/></RESULT><RESULT eventid="39" heatid="438" lane="5" points="294" resultid="3270" swimtime="00:01:17.69"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="141" birthdate="2009-01-01" firstname="Haila" gender="F" lastname="Jahn" license="423315"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="19" lane="1" points="287" resultid="141" swimtime="00:00:44.40"><SPLITS/></RESULT><RESULT eventid="9" heatid="117" lane="8" points="371" resultid="887" swimtime="00:00:32.92"><SPLITS/></RESULT><RESULT eventid="13" heatid="202" lane="7" points="309" resultid="1534" swimtime="00:01:24.95"><SPLITS><SPLIT distance="50" swimtime="00:00:40.79"/></SPLITS></RESULT><RESULT eventid="27" heatid="263" lane="5" points="315" resultid="1952" swimtime="00:00:39.62"><SPLITS/></RESULT><RESULT eventid="31" heatid="339" lane="7" points="334" resultid="2529" swimtime="00:01:32.35"><SPLITS><SPLIT distance="50" swimtime="00:00:43.70"/></SPLITS></RESULT><RESULT eventid="35" heatid="371" lane="5" points="276" resultid="2763" swimtime="00:00:37.52"><SPLITS/></RESULT><RESULT eventid="37" heatid="407" lane="1" points="329" resultid="3031" swimtime="00:02:58.65"><SPLITS><SPLIT distance="50" swimtime="00:00:41.63"/><SPLIT distance="100" swimtime="00:01:26.30"/><SPLIT distance="150" swimtime="00:02:14.54"/></SPLITS></RESULT><RESULT eventid="39" heatid="433" lane="4" points="330" resultid="3229" swimtime="00:01:14.81"><SPLITS><SPLIT distance="50" swimtime="00:00:34.69"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="143" birthdate="2008-01-01" firstname="Clara" gender="F" lastname="Welker" license="395039"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="19" lane="3" points="321" resultid="143" swimtime="00:00:42.79"><SPLITS/></RESULT><RESULT eventid="9" heatid="121" lane="5" points="378" resultid="916" swimtime="00:00:32.71"><SPLITS/></RESULT><RESULT eventid="13" heatid="200" lane="4" points="327" resultid="1515" swimtime="00:01:23.34"><SPLITS><SPLIT distance="50" swimtime="00:00:40.88"/></SPLITS></RESULT><RESULT eventid="27" heatid="266" lane="8" points="337" resultid="1979" swimtime="00:00:38.77"><SPLITS/></RESULT><RESULT eventid="29" heatid="300" lane="6" points="322" resultid="2235" swimtime="00:02:44.74"><SPLITS><SPLIT distance="50" swimtime="00:00:34.95"/><SPLIT distance="100" swimtime="00:01:17.37"/><SPLIT distance="150" swimtime="00:02:00.99"/></SPLITS></RESULT><RESULT eventid="35" heatid="374" lane="6" points="277" resultid="2788" swimtime="00:00:37.45"><SPLITS/></RESULT><RESULT eventid="39" heatid="441" lane="1" points="327" resultid="3289" swimtime="00:01:15.04"><SPLITS><SPLIT distance="50" swimtime="00:00:35.54"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="146" birthdate="2009-01-01" firstname="Mara Malin" gender="F" lastname="Walther" license="362627"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="19" lane="6" points="318" resultid="146" swimtime="00:00:42.92"><SPLITS/></RESULT><RESULT eventid="3" heatid="47" lane="4" points="360" resultid="355" swimtime="00:05:32.10"><SPLITS><SPLIT distance="100" swimtime="00:01:17.92"/><SPLIT distance="200" swimtime="00:02:42.45"/><SPLIT distance="300" swimtime="00:04:07.99"/></SPLITS></RESULT><RESULT eventid="9" heatid="120" lane="8" points="360" resultid="911" swimtime="00:00:33.26"><SPLITS/></RESULT><RESULT eventid="11" heatid="166" lane="3" points="332" resultid="1253" swimtime="00:03:02.03"><SPLITS><SPLIT distance="50" swimtime="00:00:37.49"/><SPLIT distance="100" swimtime="00:01:25.66"/><SPLIT distance="150" swimtime="00:02:22.80"/></SPLITS></RESULT><RESULT eventid="29" heatid="300" lane="5" points="362" resultid="2234" swimtime="00:02:38.44"><SPLITS><SPLIT distance="50" swimtime="00:00:36.49"/><SPLIT distance="100" swimtime="00:01:16.42"/><SPLIT distance="150" swimtime="00:01:57.62"/></SPLITS></RESULT><RESULT eventid="31" heatid="337" lane="7" points="268" resultid="2513" swimtime="00:01:39.41"><SPLITS><SPLIT distance="50" swimtime="00:00:44.94"/></SPLITS></RESULT><RESULT eventid="35" heatid="374" lane="2" points="313" resultid="2784" swimtime="00:00:35.95"><SPLITS/></RESULT><RESULT eventid="39" heatid="439" lane="2" points="355" resultid="3275" swimtime="00:01:12.97"><SPLITS><SPLIT distance="50" swimtime="00:00:35.06"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="153" birthdate="2011-01-01" firstname="Florentine" gender="F" lastname="Stein" license="450789"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="20" lane="5" points="359" resultid="153" swimtime="00:00:41.21"><SPLITS/></RESULT><RESULT eventid="7" heatid="88" lane="8" resultid="664" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="9" heatid="126" lane="3" points="494" resultid="954" swimtime="00:00:29.93"><SPLITS/></RESULT><RESULT eventid="27" heatid="269" lane="6" points="380" resultid="2000" swimtime="00:00:37.22"><SPLITS/></RESULT><RESULT eventid="29" heatid="299" lane="4" points="373" resultid="2225" swimtime="00:02:36.89"><SPLITS><SPLIT distance="50" swimtime="00:00:33.75"/><SPLIT distance="100" swimtime="00:01:12.88"/><SPLIT distance="150" swimtime="00:01:55.38"/></SPLITS></RESULT><RESULT eventid="35" heatid="377" lane="2" points="412" resultid="2807" swimtime="00:00:32.82"><SPLITS/></RESULT><RESULT eventid="39" heatid="439" lane="6" points="434" resultid="3279" swimtime="00:01:08.29"><SPLITS><SPLIT distance="50" swimtime="00:00:31.54"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="156" birthdate="2004-01-01" firstname="Julia" gender="F" lastname="Metterlein" license="357959"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="20" lane="8" points="339" resultid="156" swimtime="00:00:41.98"><SPLITS/></RESULT><RESULT eventid="9" heatid="121" lane="6" points="400" resultid="917" swimtime="00:00:32.12"><SPLITS/></RESULT><RESULT eventid="31" heatid="340" lane="6" points="362" resultid="2536" swimtime="00:01:29.94"><SPLITS><SPLIT distance="50" swimtime="00:00:42.60"/></SPLITS></RESULT><RESULT eventid="35" heatid="374" lane="1" points="282" resultid="2783" swimtime="00:00:37.23"><SPLITS/></RESULT><RESULT eventid="39" heatid="440" lane="6" points="377" resultid="3286" swimtime="00:01:11.53"><SPLITS><SPLIT distance="50" swimtime="00:00:33.93"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="157" birthdate="2001-01-01" firstname="Saskia" gender="F" lastname="Münch" license="390335"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="21" lane="1" points="261" resultid="157" swimtime="00:00:45.79"><SPLITS/></RESULT><RESULT eventid="9" heatid="122" lane="7" points="333" resultid="926" swimtime="00:00:34.12"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="167" birthdate="2003-01-01" firstname="Luana" gender="F" lastname="Liegat" license="324323"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="22" lane="4" points="451" resultid="167" swimtime="00:00:38.19"><SPLITS/></RESULT><RESULT eventid="9" heatid="127" lane="5" points="484" resultid="963" swimtime="00:00:30.14"><SPLITS/></RESULT><RESULT eventid="31" heatid="341" lane="5" points="409" resultid="2543" swimtime="00:01:26.35"><SPLITS><SPLIT distance="50" swimtime="00:00:39.77"/></SPLITS></RESULT><RESULT eventid="35" heatid="381" lane="7" points="399" resultid="2842" swimtime="00:00:33.16"><SPLITS/></RESULT><RESULT eventid="39" heatid="446" lane="7" points="450" resultid="3334" swimtime="00:01:07.46"><SPLITS><SPLIT distance="50" swimtime="00:00:31.87"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="172" birthdate="2009-01-01" firstname="Helena" gender="F" lastname="Bersch" license="383933"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="23" lane="2" points="448" resultid="172" swimtime="00:00:38.29"><SPLITS/></RESULT><RESULT eventid="7" heatid="90" lane="4" resultid="676" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="9" heatid="126" lane="1" points="400" resultid="952" swimtime="00:00:32.11"><SPLITS/></RESULT><RESULT eventid="11" heatid="172" lane="7" resultid="1305" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="29" heatid="303" lane="5" points="415" resultid="2257" swimtime="00:02:31.42"><SPLITS><SPLIT distance="50" swimtime="00:00:34.23"/><SPLIT distance="100" swimtime="00:01:12.71"/><SPLIT distance="150" swimtime="00:01:52.60"/></SPLITS></RESULT><RESULT eventid="31" heatid="343" lane="8" points="389" resultid="2562" swimtime="00:01:27.78"><SPLITS><SPLIT distance="50" swimtime="00:00:42.74"/></SPLITS></RESULT><RESULT eventid="35" heatid="379" lane="4" points="432" resultid="2823" swimtime="00:00:32.30"><SPLITS/></RESULT><RESULT eventid="39" heatid="443" lane="4" points="410" resultid="3308" swimtime="00:01:09.56"><SPLITS><SPLIT distance="50" swimtime="00:00:32.89"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="173" birthdate="2009-01-01" firstname="Helena" gender="F" lastname="Hauer" license="406750"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="23" lane="3" points="494" resultid="173" swimtime="00:00:37.05"><SPLITS/></RESULT><RESULT eventid="7" heatid="90" lane="5" points="490" resultid="677" swimtime="00:02:56.19"><SPLITS><SPLIT distance="50" swimtime="00:00:39.09"/><SPLIT distance="100" swimtime="00:01:24.14"/><SPLIT distance="150" swimtime="00:02:10.52"/></SPLITS></RESULT><RESULT eventid="9" heatid="130" lane="2" points="573" resultid="984" swimtime="00:00:28.49"><SPLITS/></RESULT><RESULT eventid="11" heatid="173" lane="7" points="530" resultid="1313" swimtime="00:02:35.78"><SPLITS><SPLIT distance="50" swimtime="00:00:33.10"/><SPLIT distance="100" swimtime="00:01:15.03"/><SPLIT distance="150" swimtime="00:02:02.20"/></SPLITS></RESULT><RESULT eventid="31" heatid="343" lane="1" points="471" resultid="2555" swimtime="00:01:22.42"><SPLITS><SPLIT distance="50" swimtime="00:00:39.17"/></SPLITS></RESULT><RESULT eventid="39" heatid="449" lane="7" points="569" resultid="3356" swimtime="00:01:02.37"><SPLITS><SPLIT distance="50" swimtime="00:00:29.59"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="175" birthdate="2000-01-01" firstname="Natalie" gender="F" lastname="Wöltinger" license="266843"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="23" lane="5" points="516" resultid="175" swimtime="00:00:36.53"><SPLITS/></RESULT><RESULT eventid="7" heatid="92" lane="5" points="601" resultid="693" swimtime="00:02:44.59"><SPLITS><SPLIT distance="50" swimtime="00:00:38.25"/><SPLIT distance="100" swimtime="00:01:20.32"/><SPLIT distance="150" swimtime="00:02:02.60"/></SPLITS></RESULT><RESULT eventid="11" heatid="174" lane="5" points="621" resultid="1319" swimtime="00:02:27.77"><SPLITS><SPLIT distance="50" swimtime="00:00:32.26"/><SPLIT distance="100" swimtime="00:01:11.65"/><SPLIT distance="150" swimtime="00:01:53.94"/></SPLITS></RESULT><RESULT eventid="15" heatid="227" lane="5" points="598" resultid="1720" swimtime="00:18:12.34"><SPLITS><SPLIT distance="100" swimtime="00:01:07.91"/><SPLIT distance="200" swimtime="00:02:19.55"/><SPLIT distance="300" swimtime="00:03:31.88"/><SPLIT distance="400" swimtime="00:04:44.18"/><SPLIT distance="500" swimtime="00:05:56.70"/><SPLIT distance="600" swimtime="00:07:09.59"/><SPLIT distance="700" swimtime="00:08:23.35"/><SPLIT distance="800" swimtime="00:09:37.36"/><SPLIT distance="900" swimtime="00:10:51.19"/><SPLIT distance="1000" swimtime="00:12:04.74"/><SPLIT distance="1100" swimtime="00:13:18.57"/><SPLIT distance="1200" swimtime="00:14:32.49"/><SPLIT distance="1300" swimtime="00:15:46.50"/><SPLIT distance="1400" swimtime="00:17:00.41"/></SPLITS></RESULT><RESULT eventid="29" heatid="307" lane="3" points="625" resultid="2285" swimtime="00:02:12.10"><SPLITS><SPLIT distance="50" swimtime="00:00:31.26"/><SPLIT distance="100" swimtime="00:01:03.74"/><SPLIT distance="150" swimtime="00:01:38.47"/></SPLITS></RESULT><RESULT eventid="31" heatid="344" lane="5" points="507" resultid="2567" swimtime="00:01:20.41"><SPLITS><SPLIT distance="50" swimtime="00:00:38.38"/></SPLITS></RESULT><RESULT eventid="41" heatid="478" lane="4" points="627" resultid="3573" swimtime="00:05:11.06"><SPLITS><SPLIT distance="50" swimtime="00:00:33.25"/><SPLIT distance="100" swimtime="00:01:11.57"/><SPLIT distance="150" swimtime="00:01:52.83"/><SPLIT distance="200" swimtime="00:02:34.24"/><SPLIT distance="250" swimtime="00:03:17.76"/><SPLIT distance="300" swimtime="00:04:01.51"/><SPLIT distance="350" swimtime="00:04:37.33"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="179" birthdate="2009-01-01" firstname="Neele" gender="F" lastname="Scharnweber" license="392894"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="24" lane="1" resultid="179" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="7" heatid="92" lane="2" resultid="690" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="9" heatid="131" lane="6" points="565" resultid="994" swimtime="00:00:28.63"><SPLITS/></RESULT><RESULT eventid="11" heatid="174" lane="2" points="591" resultid="1316" swimtime="00:02:30.27"><SPLITS><SPLIT distance="50" swimtime="00:00:32.23"/><SPLIT distance="100" swimtime="00:01:11.20"/><SPLIT distance="150" swimtime="00:01:55.24"/></SPLITS></RESULT><RESULT eventid="13" heatid="209" lane="5" points="589" resultid="1587" swimtime="00:01:08.50"><SPLITS><SPLIT distance="50" swimtime="00:00:33.27"/></SPLITS></RESULT><RESULT eventid="27" heatid="272" lane="4" points="571" resultid="2021" swimtime="00:00:32.52"><SPLITS/></RESULT><RESULT eventid="29" heatid="307" lane="7" points="580" resultid="2289" swimtime="00:02:15.44"><SPLITS><SPLIT distance="50" swimtime="00:00:31.24"/><SPLIT distance="100" swimtime="00:01:05.04"/><SPLIT distance="150" swimtime="00:01:40.63"/></SPLITS></RESULT><RESULT eventid="31" heatid="344" lane="8" points="525" resultid="2570" swimtime="00:01:19.45"><SPLITS><SPLIT distance="50" swimtime="00:00:38.16"/></SPLITS></RESULT><RESULT eventid="35" heatid="381" lane="6" points="502" resultid="2841" swimtime="00:00:30.72"><SPLITS/></RESULT><RESULT eventid="37" heatid="411" lane="6" points="574" resultid="3068" swimtime="00:02:28.38"><SPLITS><SPLIT distance="100" swimtime="00:01:11.96"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="180" birthdate="2007-01-01" firstname="Jennifer" gender="F" lastname="Thiel" license="358269"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="24" lane="2" points="466" resultid="180" swimtime="00:00:37.79"><SPLITS/></RESULT><RESULT eventid="7" heatid="92" lane="7" points="463" resultid="695" swimtime="00:02:59.61"><SPLITS><SPLIT distance="50" swimtime="00:00:39.44"/><SPLIT distance="100" swimtime="00:01:25.05"/><SPLIT distance="150" swimtime="00:02:12.06"/></SPLITS></RESULT><RESULT eventid="9" heatid="123" lane="1" resultid="928" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="31" heatid="344" lane="6" points="443" resultid="2568" swimtime="00:01:24.10"><SPLITS><SPLIT distance="50" swimtime="00:00:38.19"/></SPLITS></RESULT><RESULT eventid="39" heatid="443" lane="5" points="407" resultid="3309" swimtime="00:01:09.73"><SPLITS><SPLIT distance="50" swimtime="00:00:32.71"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="195" birthdate="2003-01-01" firstname="Josia" gender="M" lastname="Topf" license="332559"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="26" lane="6" points="63" resultid="195" swimtime="00:01:04.92"><SPLITS/></RESULT><RESULT eventid="4" heatid="53" lane="6" points="107" resultid="401" swimtime="00:07:42.58"><SPLITS><SPLIT distance="100" swimtime="00:01:49.65"/><SPLIT distance="200" swimtime="00:03:47.72"/><SPLIT distance="300" swimtime="00:05:47.25"/></SPLITS></RESULT><RESULT eventid="10" heatid="135" lane="4" points="88" resultid="1016" swimtime="00:00:46.95"><SPLITS/></RESULT><RESULT eventid="12" heatid="175" lane="2" points="98" resultid="1323" swimtime="00:04:06.91"><SPLITS><SPLIT distance="50" swimtime="00:00:54.47"/><SPLIT distance="100" swimtime="00:01:56.09"/><SPLIT distance="150" swimtime="00:03:11.39"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="198" birthdate="2016-01-01" firstname="Johannes" gender="M" lastname="Zimmermann" license="478967"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="27" lane="1" points="76" resultid="198" swimtime="00:01:01.04"><SPLITS/></RESULT><RESULT eventid="10" heatid="136" lane="6" points="116" resultid="1026" swimtime="00:00:42.82"><SPLITS/></RESULT><RESULT eventid="14" heatid="211" lane="6" points="103" resultid="1602" swimtime="00:01:50.03"><SPLITS><SPLIT distance="50" swimtime="00:00:51.58"/></SPLITS></RESULT><RESULT eventid="28" heatid="276" lane="7" points="106" resultid="2053" swimtime="00:00:49.99"><SPLITS/></RESULT><RESULT eventid="30" heatid="310" lane="5" points="91" resultid="2308" swimtime="00:03:46.46"><SPLITS><SPLIT distance="50" swimtime="00:00:48.18"/><SPLIT distance="100" swimtime="00:01:46.35"/><SPLIT distance="150" swimtime="00:02:47.32"/></SPLITS></RESULT><RESULT eventid="36" heatid="384" lane="7" points="51" resultid="2861" swimtime="00:01:00.00"><SPLITS/></RESULT><RESULT eventid="38" heatid="413" lane="3" points="114" resultid="3079" swimtime="00:03:50.72"><SPLITS><SPLIT distance="50" swimtime="00:00:53.43"/><SPLIT distance="100" swimtime="00:01:53.31"/><SPLIT distance="150" swimtime="00:02:54.87"/></SPLITS></RESULT><RESULT eventid="40" heatid="454" lane="6" points="93" resultid="3395" swimtime="00:01:43.36"><SPLITS><SPLIT distance="50" swimtime="00:00:47.95"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="199" birthdate="2015-01-01" firstname="Jonathan" gender="M" lastname="Jakubietz" license="475247"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="27" lane="2" points="79" resultid="199" swimtime="00:01:00.30"><SPLITS/></RESULT><RESULT eventid="10" heatid="136" lane="4" points="129" resultid="1024" swimtime="00:00:41.28"><SPLITS/></RESULT><RESULT eventid="14" heatid="212" lane="8" points="97" resultid="1612" swimtime="00:01:52.16"><SPLITS><SPLIT distance="50" swimtime="00:00:54.46"/></SPLITS></RESULT><RESULT eventid="28" heatid="275" lane="4" points="112" resultid="2042" swimtime="00:00:49.17"><SPLITS/></RESULT><RESULT eventid="30" heatid="310" lane="8" points="79" resultid="2311" swimtime="00:03:57.16"><SPLITS><SPLIT distance="50" swimtime="00:00:50.38"/><SPLIT distance="100" swimtime="00:01:51.16"/><SPLIT distance="150" swimtime="00:02:57.72"/></SPLITS></RESULT><RESULT eventid="36" heatid="383" lane="5" points="48" resultid="2854" swimtime="00:01:00.93"><SPLITS/></RESULT><RESULT eventid="40" heatid="454" lane="8" points="82" resultid="3397" swimtime="00:01:47.67"><SPLITS><SPLIT distance="50" swimtime="00:00:49.40"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="207" birthdate="2012-01-01" firstname="Constantin" gender="M" lastname="Jakubietz" license="446968"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="28" lane="3" points="103" resultid="207" swimtime="00:00:55.21"><SPLITS/></RESULT><RESULT eventid="10" heatid="139" lane="4" points="182" resultid="1047" swimtime="00:00:36.86"><SPLITS/></RESULT><RESULT eventid="14" heatid="214" lane="4" points="145" resultid="1624" swimtime="00:01:38.02"><SPLITS><SPLIT distance="50" swimtime="00:00:46.30"/></SPLITS></RESULT><RESULT eventid="28" heatid="279" lane="8" resultid="2076" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="36" heatid="386" lane="1" resultid="2871" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="40" heatid="456" lane="4" resultid="3409" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="210" birthdate="2014-01-01" firstname="Florian" gender="M" lastname="Wegner" license="460206"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="28" lane="6" points="102" resultid="210" swimtime="00:00:55.38"><SPLITS/></RESULT><RESULT eventid="10" heatid="136" lane="3" points="123" resultid="1023" swimtime="00:00:42.02"><SPLITS/></RESULT><RESULT eventid="14" heatid="212" lane="2" points="110" resultid="1606" swimtime="00:01:47.64"><SPLITS><SPLIT distance="50" swimtime="00:00:51.75"/></SPLITS></RESULT><RESULT eventid="28" heatid="277" lane="2" points="119" resultid="2055" swimtime="00:00:48.12"><SPLITS/></RESULT><RESULT eventid="32" heatid="346" lane="3" points="97" resultid="2577" swimtime="00:02:03.40"><SPLITS><SPLIT distance="50" swimtime="00:00:59.42"/></SPLITS></RESULT><RESULT eventid="40" heatid="455" lane="8" points="116" resultid="3405" swimtime="00:01:35.82"><SPLITS><SPLIT distance="50" swimtime="00:00:48.01"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="211" birthdate="2013-01-01" firstname="Rémi" gender="M" lastname="Lahner" license="460138"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="28" lane="7" points="82" resultid="211" swimtime="00:00:59.63"><SPLITS/></RESULT><RESULT eventid="10" heatid="136" lane="2" points="110" resultid="1022" swimtime="00:00:43.64"><SPLITS/></RESULT><RESULT eventid="14" heatid="211" lane="3" points="110" resultid="1600" swimtime="00:01:47.40"><SPLITS><SPLIT distance="50" swimtime="00:00:49.96"/></SPLITS></RESULT><RESULT eventid="28" heatid="276" lane="3" points="109" resultid="2049" swimtime="00:00:49.56"><SPLITS/></RESULT><RESULT eventid="40" heatid="454" lane="2" points="121" resultid="3391" swimtime="00:01:34.59"><SPLITS><SPLIT distance="50" swimtime="00:00:44.74"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="217" birthdate="2013-01-01" firstname="Philipp" gender="M" lastname="Böhm" license="460131"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="29" lane="5" resultid="217" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="10" heatid="138" lane="2" resultid="1038" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="14" heatid="214" lane="8" resultid="1628" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="224" birthdate="2014-01-01" firstname="Fedor" gender="M" lastname="Mikhalenko" license="474609"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="30" lane="4" points="128" resultid="224" swimtime="00:00:51.47"><SPLITS/></RESULT><RESULT comment="12:38 Start vor dem Startsignal" eventid="8" heatid="94" lane="4" resultid="707" status="DSQ" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="10" heatid="139" lane="3" points="139" resultid="1046" swimtime="00:00:40.29"><SPLITS/></RESULT><RESULT eventid="12" heatid="176" lane="3" points="169" resultid="1330" swimtime="00:03:25.87"><SPLITS><SPLIT distance="50" swimtime="00:00:52.62"/><SPLIT distance="100" swimtime="00:01:42.09"/><SPLIT distance="150" swimtime="00:02:42.20"/></SPLITS></RESULT><RESULT eventid="28" heatid="279" lane="6" points="149" resultid="2074" swimtime="00:00:44.69"><SPLITS/></RESULT><RESULT eventid="32" heatid="348" lane="5" points="132" resultid="2594" swimtime="00:01:51.68"><SPLITS><SPLIT distance="50" swimtime="00:00:53.46"/></SPLITS></RESULT><RESULT eventid="38" heatid="415" lane="4" points="204" resultid="3094" swimtime="00:03:09.93"><SPLITS><SPLIT distance="50" swimtime="00:00:45.83"/><SPLIT distance="100" swimtime="00:01:34.79"/><SPLIT distance="150" swimtime="00:02:23.63"/></SPLITS></RESULT><RESULT eventid="40" heatid="455" lane="4" points="175" resultid="3401" swimtime="00:01:23.72"><SPLITS><SPLIT distance="50" swimtime="00:00:40.76"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="228" birthdate="2010-01-01" firstname="Mateo" gender="M" lastname="Gärtner" license="473812"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="30" lane="8" resultid="228" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="8" heatid="94" lane="3" points="156" resultid="706" swimtime="00:03:53.94"><SPLITS><SPLIT distance="50" swimtime="00:00:52.46"/><SPLIT distance="100" swimtime="00:01:52.92"/><SPLIT distance="150" swimtime="00:02:57.17"/></SPLITS></RESULT><RESULT eventid="10" heatid="142" lane="1" points="194" resultid="1067" swimtime="00:00:36.12"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="234" birthdate="2015-01-01" firstname="Paul" gender="M" lastname="Holzinger" license="474974"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="31" lane="6" points="133" resultid="234" swimtime="00:00:50.78"><SPLITS/></RESULT><RESULT eventid="4" heatid="55" lane="8" points="164" resultid="417" swimtime="00:06:41.81"><SPLITS><SPLIT distance="100" swimtime="00:01:37.21"/><SPLIT distance="200" swimtime="00:03:22.50"/><SPLIT distance="300" swimtime="00:05:06.00"/></SPLITS></RESULT><RESULT eventid="10" heatid="138" lane="3" points="150" resultid="1039" swimtime="00:00:39.30"><SPLITS/></RESULT><RESULT eventid="12" heatid="175" lane="4" points="151" resultid="1325" swimtime="00:03:33.76"><SPLITS><SPLIT distance="50" swimtime="00:00:48.00"/><SPLIT distance="100" swimtime="00:01:44.98"/><SPLIT distance="150" swimtime="00:02:47.01"/></SPLITS></RESULT><RESULT eventid="30" heatid="312" lane="5" points="159" resultid="2323" swimtime="00:03:08.03"><SPLITS><SPLIT distance="50" swimtime="00:00:45.91"/><SPLIT distance="100" swimtime="00:01:35.27"/><SPLIT distance="150" swimtime="00:02:24.73"/></SPLITS></RESULT><RESULT eventid="36" heatid="386" lane="4" points="107" resultid="2874" swimtime="00:00:46.78"><SPLITS/></RESULT><RESULT eventid="40" heatid="457" lane="2" points="153" resultid="3414" swimtime="00:01:27.55"><SPLITS><SPLIT distance="50" swimtime="00:00:44.23"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="235" birthdate="2013-01-01" firstname="Thadeo" gender="M" lastname="Puchalla" license="475933"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="31" lane="7" points="134" resultid="235" swimtime="00:00:50.67"><SPLITS/></RESULT><RESULT eventid="10" heatid="139" lane="1" points="126" resultid="1044" swimtime="00:00:41.62"><SPLITS/></RESULT><RESULT eventid="14" heatid="211" lane="7" points="113" resultid="1603" swimtime="00:01:46.43"><SPLITS><SPLIT distance="50" swimtime="00:00:49.93"/></SPLITS></RESULT><RESULT eventid="28" heatid="276" lane="1" points="120" resultid="2047" swimtime="00:00:47.98"><SPLITS/></RESULT><RESULT eventid="30" heatid="310" lane="7" points="101" resultid="2310" swimtime="00:03:38.75"><SPLITS><SPLIT distance="50" swimtime="00:00:47.73"/><SPLIT distance="100" swimtime="00:01:45.56"/><SPLIT distance="150" swimtime="00:02:45.71"/></SPLITS></RESULT><RESULT eventid="32" heatid="347" lane="6" points="150" resultid="2587" swimtime="00:01:46.86"><SPLITS><SPLIT distance="50" swimtime="00:00:51.23"/></SPLITS></RESULT><RESULT eventid="36" heatid="383" lane="4" points="87" resultid="2853" swimtime="00:00:50.16"><SPLITS/></RESULT><RESULT eventid="40" heatid="455" lane="2" points="121" resultid="3399" swimtime="00:01:34.69"><SPLITS><SPLIT distance="50" swimtime="00:00:44.73"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="237" birthdate="2008-01-01" firstname="Rene" gender="M" lastname="Thiel" license="389089"><HANDICAP/><ENTRIES/><RESULTS><RESULT comment="09:44 Start vor dem Startsginal" eventid="2" heatid="32" lane="1" resultid="237" status="DSQ" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="10" heatid="143" lane="5" points="363" resultid="1078" swimtime="00:00:29.30"><SPLITS/></RESULT><RESULT eventid="30" heatid="317" lane="2" points="314" resultid="2359" swimtime="00:02:29.97"><SPLITS><SPLIT distance="50" swimtime="00:00:30.95"/><SPLIT distance="100" swimtime="00:01:08.55"/><SPLIT distance="150" swimtime="00:01:50.46"/></SPLITS></RESULT><RESULT eventid="36" heatid="387" lane="5" points="335" resultid="2882" swimtime="00:00:32.06"><SPLITS/></RESULT><RESULT eventid="40" heatid="460" lane="7" points="395" resultid="3442" swimtime="00:01:03.82"><SPLITS><SPLIT distance="50" swimtime="00:00:29.87"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="240" birthdate="2012-01-01" firstname="Julius" gender="M" lastname="Wöhler" license="446973"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="32" lane="4" resultid="240" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="4" heatid="57" lane="6" resultid="431" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="10" heatid="143" lane="2" resultid="1075" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="12" heatid="177" lane="2" resultid="1337" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="241" birthdate="2010-01-01" firstname="Julian" gender="M" lastname="Jakubietz" license="447010"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="32" lane="5" points="210" resultid="241" swimtime="00:00:43.62"><SPLITS/></RESULT><RESULT eventid="10" heatid="146" lane="3" points="315" resultid="1100" swimtime="00:00:30.70"><SPLITS/></RESULT><RESULT eventid="12" heatid="180" lane="5" points="268" resultid="1362" swimtime="00:02:56.75"><SPLITS><SPLIT distance="50" swimtime="00:00:38.49"/><SPLIT distance="100" swimtime="00:01:23.47"/><SPLIT distance="150" swimtime="00:02:18.60"/></SPLITS></RESULT><RESULT eventid="30" heatid="319" lane="6" points="296" resultid="2379" swimtime="00:02:33.03"><SPLITS><SPLIT distance="50" swimtime="00:00:34.26"/><SPLIT distance="100" swimtime="00:01:13.50"/><SPLIT distance="150" swimtime="00:01:55.40"/></SPLITS></RESULT><RESULT eventid="36" heatid="389" lane="4" points="240" resultid="2897" swimtime="00:00:35.82"><SPLITS/></RESULT><RESULT eventid="40" heatid="466" lane="1" points="320" resultid="3483" swimtime="00:01:08.46"><SPLITS><SPLIT distance="50" swimtime="00:00:33.03"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="248" birthdate="2010-01-01" firstname="Andreas" gender="M" lastname="Wegner" license="438077"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="33" lane="4" points="235" resultid="248" swimtime="00:00:42.01"><SPLITS/></RESULT><RESULT eventid="6" heatid="74" lane="2" points="181" resultid="552" swimtime="00:01:27.32"><SPLITS><SPLIT distance="50" swimtime="00:00:40.83"/></SPLITS></RESULT><RESULT eventid="10" heatid="146" lane="8" points="278" resultid="1105" swimtime="00:00:32.02"><SPLITS/></RESULT><RESULT eventid="28" heatid="283" lane="8" points="218" resultid="2108" swimtime="00:00:39.37"><SPLITS/></RESULT><RESULT eventid="30" heatid="318" lane="1" points="255" resultid="2366" swimtime="00:02:40.66"><SPLITS><SPLIT distance="50" swimtime="00:00:37.41"/><SPLIT distance="100" swimtime="00:01:18.07"/><SPLIT distance="150" swimtime="00:02:01.04"/></SPLITS></RESULT><RESULT eventid="36" heatid="391" lane="6" points="204" resultid="2915" swimtime="00:00:37.78"><SPLITS/></RESULT><RESULT eventid="40" heatid="459" lane="4" points="285" resultid="3432" swimtime="00:01:11.16"><SPLITS><SPLIT distance="50" swimtime="00:00:35.02"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="249" birthdate="2013-01-01" firstname="Filip" gender="M" lastname="Lazic" license="470933"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="33" lane="5" points="212" resultid="249" swimtime="00:00:43.52"><SPLITS/></RESULT><RESULT eventid="8" heatid="96" lane="5" points="237" resultid="722" swimtime="00:03:23.49"><SPLITS><SPLIT distance="50" swimtime="00:00:46.03"/><SPLIT distance="100" swimtime="00:01:38.35"/><SPLIT distance="150" swimtime="00:02:31.28"/></SPLITS></RESULT><RESULT eventid="12" heatid="179" lane="6" points="224" resultid="1355" swimtime="00:03:07.61"><SPLITS><SPLIT distance="50" swimtime="00:00:45.85"/><SPLIT distance="100" swimtime="00:01:32.36"/><SPLIT distance="150" swimtime="00:02:25.42"/></SPLITS></RESULT><RESULT eventid="14" heatid="216" lane="2" points="207" resultid="1636" swimtime="00:01:27.15"><SPLITS><SPLIT distance="50" swimtime="00:00:43.55"/></SPLITS></RESULT><RESULT eventid="28" heatid="281" lane="8" points="209" resultid="2092" swimtime="00:00:39.90"><SPLITS/></RESULT><RESULT eventid="30" heatid="314" lane="8" points="205" resultid="2341" swimtime="00:02:52.79"><SPLITS><SPLIT distance="50" swimtime="00:00:39.22"/><SPLIT distance="100" swimtime="00:01:22.77"/><SPLIT distance="150" swimtime="00:02:09.87"/></SPLITS></RESULT><RESULT eventid="38" heatid="416" lane="1" points="232" resultid="3099" swimtime="00:03:01.96"><SPLITS><SPLIT distance="50" swimtime="00:00:44.55"/><SPLIT distance="100" swimtime="00:01:30.36"/><SPLIT distance="150" swimtime="00:02:18.40"/></SPLITS></RESULT><RESULT eventid="40" heatid="461" lane="4" points="201" resultid="3447" swimtime="00:01:19.91"><SPLITS><SPLIT distance="50" swimtime="00:00:38.24"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="256" birthdate="2011-01-01" firstname="Ivan" gender="M" lastname="Vasylyna" license="453314"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="34" lane="4" points="199" resultid="256" swimtime="00:00:44.40"><SPLITS/></RESULT><RESULT eventid="8" heatid="97" lane="7" points="226" resultid="732" swimtime="00:03:26.50"><SPLITS><SPLIT distance="50" swimtime="00:00:46.67"/><SPLIT distance="100" swimtime="00:01:41.29"/><SPLIT distance="150" swimtime="00:02:34.15"/></SPLITS></RESULT><RESULT eventid="10" heatid="145" lane="1" points="266" resultid="1090" swimtime="00:00:32.49"><SPLITS/></RESULT><RESULT eventid="12" heatid="180" lane="2" points="250" resultid="1359" swimtime="00:03:00.77"><SPLITS><SPLIT distance="50" swimtime="00:00:42.46"/><SPLIT distance="100" swimtime="00:01:27.07"/><SPLIT distance="150" swimtime="00:02:21.52"/></SPLITS></RESULT><RESULT eventid="28" heatid="281" lane="7" points="218" resultid="2091" swimtime="00:00:39.39"><SPLITS/></RESULT><RESULT eventid="30" heatid="321" lane="8" points="271" resultid="2395" swimtime="00:02:37.49"><SPLITS><SPLIT distance="50" swimtime="00:00:37.01"/><SPLIT distance="100" swimtime="00:01:17.02"/><SPLIT distance="150" swimtime="00:01:59.57"/></SPLITS></RESULT><RESULT eventid="32" heatid="351" lane="8" points="191" resultid="2619" swimtime="00:01:38.71"><SPLITS><SPLIT distance="50" swimtime="00:00:47.76"/></SPLITS></RESULT><RESULT comment="14:28 Der Sportler brachte mehrfach die Arme nicht gleichzeitig nach vorne" eventid="36" heatid="387" lane="6" resultid="2883" status="DSQ" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="40" heatid="464" lane="1" points="253" resultid="3467" swimtime="00:01:14.07"><SPLITS><SPLIT distance="50" swimtime="00:00:36.55"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="259" birthdate="2012-01-01" firstname="Amir" gender="M" lastname="Gadhgadhi" license="447238"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="35" lane="1" points="203" resultid="259" swimtime="00:00:44.14"><SPLITS/></RESULT><RESULT eventid="8" heatid="96" lane="7" points="198" resultid="724" swimtime="00:03:36.00"><SPLITS><SPLIT distance="50" swimtime="00:00:45.32"/><SPLIT distance="100" swimtime="00:01:42.28"/><SPLIT distance="150" swimtime="00:02:39.31"/></SPLITS></RESULT><RESULT eventid="10" heatid="144" lane="4" points="221" resultid="1085" swimtime="00:00:34.56"><SPLITS/></RESULT><RESULT eventid="14" heatid="219" lane="1" points="163" resultid="1659" swimtime="00:01:34.43"><SPLITS><SPLIT distance="50" swimtime="00:00:45.34"/></SPLITS></RESULT><RESULT eventid="28" heatid="281" lane="4" points="200" resultid="2088" swimtime="00:00:40.53"><SPLITS/></RESULT><RESULT eventid="30" heatid="318" lane="7" points="215" resultid="2372" swimtime="00:02:50.05"><SPLITS><SPLIT distance="50" swimtime="00:00:35.82"/><SPLIT distance="100" swimtime="00:01:19.77"/><SPLIT distance="150" swimtime="00:02:06.09"/></SPLITS></RESULT><RESULT eventid="32" heatid="350" lane="7" points="183" resultid="2610" swimtime="00:01:40.02"><SPLITS><SPLIT distance="50" swimtime="00:00:46.54"/></SPLITS></RESULT><RESULT eventid="40" heatid="463" lane="7" points="205" resultid="3465" swimtime="00:01:19.42"><SPLITS><SPLIT distance="50" swimtime="00:00:36.64"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="278" birthdate="2011-01-01" firstname="Anton" gender="M" lastname="Cao" license="417199"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="37" lane="4" resultid="278" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="8" heatid="100" lane="4" resultid="752" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="12" heatid="186" lane="3" resultid="1406" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="14" heatid="222" lane="6" resultid="1687" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="30" heatid="320" lane="2" resultid="2383" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="32" heatid="354" lane="3" resultid="2637" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="38" heatid="418" lane="2" resultid="3115" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="42" heatid="480" lane="2" resultid="3586" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="280" birthdate="2005-01-01" firstname="Julian" gender="M" lastname="van Geemert" license="409353"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="37" lane="6" points="312" resultid="280" swimtime="00:00:38.25"><SPLITS/></RESULT><RESULT eventid="6" heatid="77" lane="6" points="299" resultid="580" swimtime="00:01:13.94"><SPLITS><SPLIT distance="50" swimtime="00:00:31.92"/></SPLITS></RESULT><RESULT eventid="10" heatid="151" lane="4" points="430" resultid="1141" swimtime="00:00:27.69"><SPLITS/></RESULT><RESULT eventid="12" heatid="186" lane="7" points="361" resultid="1410" swimtime="00:02:39.99"><SPLITS><SPLIT distance="50" swimtime="00:00:31.61"/><SPLIT distance="100" swimtime="00:01:14.99"/><SPLIT distance="150" swimtime="00:02:01.84"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="284" birthdate="2006-01-01" firstname="Alexander" gender="M" lastname="Primorac" license="392226"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="38" lane="2" points="428" resultid="284" swimtime="00:00:34.43"><SPLITS/></RESULT><RESULT eventid="6" heatid="77" lane="1" points="389" resultid="575" swimtime="00:01:07.72"><SPLITS><SPLIT distance="50" swimtime="00:00:31.80"/></SPLITS></RESULT><RESULT eventid="10" heatid="156" lane="6" points="517" resultid="1181" swimtime="00:00:26.04"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="289" birthdate="2008-01-01" firstname="Justus" gender="M" lastname="Lemle" license="389520"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="38" lane="7" points="391" resultid="289" swimtime="00:00:35.47"><SPLITS/></RESULT><RESULT eventid="6" heatid="74" lane="7" points="208" resultid="557" swimtime="00:01:23.40"><SPLITS><SPLIT distance="50" swimtime="00:00:36.35"/></SPLITS></RESULT><RESULT eventid="10" heatid="149" lane="3" points="350" resultid="1124" swimtime="00:00:29.65"><SPLITS/></RESULT><RESULT eventid="12" heatid="185" lane="4" points="302" resultid="1399" swimtime="00:02:49.73"><SPLITS><SPLIT distance="50" swimtime="00:00:34.57"/><SPLIT distance="100" swimtime="00:01:22.90"/><SPLIT distance="150" swimtime="00:02:09.78"/></SPLITS></RESULT><RESULT eventid="32" heatid="354" lane="6" points="345" resultid="2640" swimtime="00:01:21.04"><SPLITS><SPLIT distance="50" swimtime="00:00:38.17"/></SPLITS></RESULT><RESULT eventid="36" heatid="393" lane="3" points="297" resultid="2928" swimtime="00:00:33.36"><SPLITS/></RESULT><RESULT eventid="40" heatid="468" lane="1" points="332" resultid="3498" swimtime="00:01:07.62"><SPLITS><SPLIT distance="50" swimtime="00:00:32.35"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="292" birthdate="2007-01-01" firstname="Ben Clement" gender="M" lastname="Ying" license="372887"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="39" lane="2" points="485" resultid="292" swimtime="00:00:33.01"><SPLITS/></RESULT><RESULT eventid="10" heatid="154" lane="1" points="461" resultid="1162" swimtime="00:00:27.06"><SPLITS/></RESULT><RESULT eventid="28" heatid="287" lane="2" points="538" resultid="2133" swimtime="00:00:29.15"><SPLITS/></RESULT><RESULT eventid="36" heatid="398" lane="2" points="491" resultid="2967" swimtime="00:00:28.22"><SPLITS/></RESULT><RESULT eventid="40" heatid="472" lane="3" points="514" resultid="3532" swimtime="00:00:58.47"><SPLITS><SPLIT distance="50" swimtime="00:00:28.05"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="293" birthdate="2003-01-01" firstname="Jan" gender="M" lastname="Sedlacek" license="315494"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="39" lane="3" points="446" resultid="293" swimtime="00:00:33.96"><SPLITS/></RESULT><RESULT eventid="10" heatid="152" lane="3" resultid="1148" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="14" heatid="223" lane="5" resultid="1694" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="28" heatid="285" lane="3" resultid="2118" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="36" heatid="398" lane="3" resultid="2968" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="38" heatid="418" lane="4" resultid="3117" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="300" birthdate="2000-01-01" firstname="Eric" gender="M" lastname="Martin" license="299708"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="40" lane="2" points="519" resultid="300" swimtime="00:00:32.29"><SPLITS/></RESULT><RESULT eventid="6" heatid="78" lane="6" points="369" resultid="587" swimtime="00:01:08.94"><SPLITS><SPLIT distance="50" swimtime="00:00:28.61"/></SPLITS></RESULT><RESULT eventid="10" heatid="155" lane="6" points="499" resultid="1173" swimtime="00:00:26.35"><SPLITS/></RESULT><RESULT eventid="32" heatid="356" lane="8" points="461" resultid="2657" swimtime="00:01:13.58"><SPLITS><SPLIT distance="50" swimtime="00:00:33.27"/></SPLITS></RESULT><RESULT eventid="36" heatid="399" lane="7" points="512" resultid="2980" swimtime="00:00:27.83"><SPLITS/></RESULT><RESULT eventid="40" heatid="473" lane="3" points="510" resultid="3539" swimtime="00:00:58.64"><SPLITS><SPLIT distance="50" swimtime="00:00:27.88"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="301" birthdate="2002-01-01" firstname="Valentin" gender="M" lastname="Schmiedel" license="289162"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="40" lane="3" points="574" resultid="301" swimtime="00:00:31.21"><SPLITS/></RESULT><RESULT eventid="8" heatid="101" lane="2" points="498" resultid="758" swimtime="00:02:38.84"><SPLITS><SPLIT distance="50" swimtime="00:00:34.83"/><SPLIT distance="100" swimtime="00:01:15.05"/><SPLIT distance="150" swimtime="00:01:57.58"/></SPLITS></RESULT><RESULT eventid="10" heatid="152" lane="1" points="425" resultid="1146" swimtime="00:00:27.80"><SPLITS/></RESULT><RESULT eventid="12" heatid="189" lane="8" points="418" resultid="1434" swimtime="00:02:32.46"><SPLITS><SPLIT distance="50" swimtime="00:00:31.31"/><SPLIT distance="100" swimtime="00:01:14.05"/><SPLIT distance="150" swimtime="00:01:56.03"/></SPLITS></RESULT><RESULT eventid="32" heatid="356" lane="6" points="498" resultid="2655" swimtime="00:01:11.76"><SPLITS><SPLIT distance="50" swimtime="00:00:33.27"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="303" birthdate="2007-01-01" firstname="Magnus" gender="M" lastname="Lemle" license="372889"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="40" lane="5" points="517" resultid="303" swimtime="00:00:32.33"><SPLITS/></RESULT><RESULT eventid="8" heatid="101" lane="4" points="509" resultid="760" swimtime="00:02:37.71"><SPLITS><SPLIT distance="50" swimtime="00:00:35.66"/><SPLIT distance="100" swimtime="00:01:15.17"/><SPLIT distance="150" swimtime="00:01:56.08"/></SPLITS></RESULT><RESULT eventid="10" heatid="154" lane="2" points="463" resultid="1163" swimtime="00:00:27.02"><SPLITS/></RESULT><RESULT eventid="12" heatid="189" lane="3" points="483" resultid="1430" swimtime="00:02:25.23"><SPLITS><SPLIT distance="50" swimtime="00:00:31.13"/><SPLIT distance="100" swimtime="00:01:09.64"/><SPLIT distance="150" swimtime="00:01:51.99"/></SPLITS></RESULT><RESULT eventid="28" heatid="286" lane="3" points="409" resultid="2126" swimtime="00:00:31.92"><SPLITS/></RESULT><RESULT eventid="32" heatid="356" lane="4" points="484" resultid="2653" swimtime="00:01:12.42"><SPLITS><SPLIT distance="50" swimtime="00:00:33.56"/></SPLITS></RESULT><RESULT eventid="38" heatid="419" lane="6" points="447" resultid="3124" swimtime="00:02:26.31"><SPLITS><SPLIT distance="50" swimtime="00:00:33.77"/><SPLIT distance="100" swimtime="00:01:11.40"/><SPLIT distance="150" swimtime="00:01:49.00"/></SPLITS></RESULT><RESULT eventid="42" heatid="481" lane="5" points="516" resultid="3594" swimtime="00:05:04.01"><SPLITS><SPLIT distance="50" swimtime="00:00:31.67"/><SPLIT distance="100" swimtime="00:01:10.12"/><SPLIT distance="150" swimtime="00:01:51.52"/><SPLIT distance="200" swimtime="00:02:31.08"/><SPLIT distance="250" swimtime="00:03:13.51"/><SPLIT distance="300" swimtime="00:03:55.44"/><SPLIT distance="350" swimtime="00:04:30.51"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="311" birthdate="2014-01-01" firstname="Helena" gender="F" lastname="Gold" license="479146"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="42" lane="1" points="235" resultid="312" swimtime="00:06:22.88"><SPLITS><SPLIT distance="100" swimtime="00:01:30.69"/><SPLIT distance="200" swimtime="00:03:09.50"/><SPLIT distance="300" swimtime="00:04:48.40"/></SPLITS></RESULT><RESULT eventid="9" heatid="112" lane="7" points="243" resultid="847" swimtime="00:00:37.88"><SPLITS/></RESULT><RESULT eventid="13" heatid="197" lane="4" points="210" resultid="1491" swimtime="00:01:36.57"><SPLITS><SPLIT distance="50" swimtime="00:00:46.96"/></SPLITS></RESULT><RESULT eventid="27" heatid="260" lane="5" points="210" resultid="1928" swimtime="00:00:45.34"><SPLITS/></RESULT><RESULT eventid="29" heatid="291" lane="3" points="229" resultid="2160" swimtime="00:03:04.63"><SPLITS><SPLIT distance="50" swimtime="00:00:42.54"/><SPLIT distance="100" swimtime="00:01:30.08"/><SPLIT distance="150" swimtime="00:02:18.47"/></SPLITS></RESULT><RESULT eventid="35" heatid="365" lane="1" points="110" resultid="2711" swimtime="00:00:50.97"><SPLITS/></RESULT><RESULT eventid="37" heatid="404" lane="6" points="242" resultid="3012" swimtime="00:03:17.76"><SPLITS><SPLIT distance="50" swimtime="00:00:48.47"/><SPLIT distance="100" swimtime="00:01:39.26"/><SPLIT distance="150" swimtime="00:02:29.86"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="329" birthdate="2014-01-01" firstname="Pauline" gender="F" lastname="Ziegler" license="470932"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="44" lane="8" points="296" resultid="335" swimtime="00:05:54.46"><SPLITS><SPLIT distance="100" swimtime="00:01:22.08"/><SPLIT distance="200" swimtime="00:02:52.68"/><SPLIT distance="300" swimtime="00:04:25.58"/></SPLITS></RESULT><RESULT eventid="9" heatid="115" lane="5" points="285" resultid="869" swimtime="00:00:35.96"><SPLITS/></RESULT><RESULT comment="15:15 Die Teilstrecke Brust wurde nicht mit beiden Händen gleichzeitig beendet" eventid="11" heatid="160" lane="8" resultid="1210" status="DSQ" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="29" heatid="295" lane="5" points="312" resultid="2194" swimtime="00:02:46.47"><SPLITS><SPLIT distance="50" swimtime="00:00:38.84"/><SPLIT distance="100" swimtime="00:01:22.27"/><SPLIT distance="150" swimtime="00:02:06.03"/></SPLITS></RESULT><RESULT eventid="35" heatid="366" lane="4" points="129" resultid="2722" swimtime="00:00:48.30"><SPLITS/></RESULT><RESULT eventid="39" heatid="434" lane="6" points="299" resultid="3239" swimtime="00:01:17.29"><SPLITS><SPLIT distance="50" swimtime="00:00:36.52"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="336" birthdate="2011-01-01" firstname="Augusta Sofia" gender="F" lastname="Baker-Duly" license="436698"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="46" lane="2" resultid="345" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="9" heatid="121" lane="3" resultid="914" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="11" heatid="165" lane="4" resultid="1246" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="13" heatid="201" lane="6" resultid="1525" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="27" heatid="265" lane="7" resultid="1970" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="35" heatid="374" lane="3" resultid="2785" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="39" heatid="440" lane="8" resultid="3288" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="338" birthdate="2013-01-01" firstname="Ida" gender="F" lastname="Finke" license="446399"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="46" lane="5" points="285" resultid="348" swimtime="00:05:59.22"><SPLITS><SPLIT distance="100" swimtime="00:01:21.65"/><SPLIT distance="200" swimtime="00:02:55.32"/><SPLIT distance="300" swimtime="00:04:29.60"/></SPLITS></RESULT><RESULT eventid="9" heatid="122" lane="5" points="419" resultid="924" swimtime="00:00:31.62"><SPLITS/></RESULT><RESULT eventid="11" heatid="166" lane="5" points="311" resultid="1255" swimtime="00:03:06.10"><SPLITS><SPLIT distance="50" swimtime="00:00:39.15"/><SPLIT distance="100" swimtime="00:01:26.84"/><SPLIT distance="150" swimtime="00:02:25.42"/></SPLITS></RESULT><RESULT eventid="23" heatid="243" lane="4" resultid="1810" swimtime="00:00:47.56"><SPLITS/></RESULT><RESULT eventid="29" heatid="301" lane="5" points="311" resultid="2241" swimtime="00:02:46.62"><SPLITS><SPLIT distance="50" swimtime="00:00:35.51"/><SPLIT distance="100" swimtime="00:01:17.76"/><SPLIT distance="150" swimtime="00:02:03.37"/></SPLITS></RESULT><RESULT eventid="35" heatid="373" lane="4" points="310" resultid="2778" swimtime="00:00:36.07"><SPLITS/></RESULT><RESULT eventid="39" heatid="440" lane="4" points="387" resultid="3284" swimtime="00:01:10.90"><SPLITS><SPLIT distance="50" swimtime="00:00:32.75"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="346" birthdate="2010-01-01" firstname="Sophie" gender="F" lastname="Böller" license="420812"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="48" lane="5" points="349" resultid="363" swimtime="00:05:35.69"><SPLITS><SPLIT distance="100" swimtime="00:01:17.57"/><SPLIT distance="200" swimtime="00:02:42.29"/><SPLIT distance="300" swimtime="00:04:09.76"/></SPLITS></RESULT><RESULT eventid="9" heatid="127" lane="4" points="512" resultid="962" swimtime="00:00:29.58"><SPLITS/></RESULT><RESULT eventid="13" heatid="205" lane="1" points="385" resultid="1552" swimtime="00:01:18.95"><SPLITS><SPLIT distance="50" swimtime="00:00:38.16"/></SPLITS></RESULT><RESULT eventid="27" heatid="271" lane="6" points="417" resultid="2015" swimtime="00:00:36.11"><SPLITS/></RESULT><RESULT eventid="31" heatid="339" lane="6" points="337" resultid="2528" swimtime="00:01:32.14"><SPLITS><SPLIT distance="50" swimtime="00:00:43.35"/></SPLITS></RESULT><RESULT eventid="35" heatid="378" lane="1" points="393" resultid="2812" swimtime="00:00:33.35"><SPLITS/></RESULT><RESULT eventid="37" heatid="411" lane="2" points="381" resultid="3064" swimtime="00:02:50.02"><SPLITS><SPLIT distance="100" swimtime="00:01:21.55"/></SPLITS></RESULT><RESULT eventid="39" heatid="442" lane="3" points="414" resultid="3299" swimtime="00:01:09.38"><SPLITS><SPLIT distance="50" swimtime="00:00:32.77"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="350" birthdate="2013-01-01" firstname="Coralie-Sophie" gender="F" lastname="Walther" license="425763"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="49" lane="1" points="398" resultid="367" swimtime="00:05:21.32"><SPLITS><SPLIT distance="100" swimtime="00:01:15.00"/><SPLIT distance="200" swimtime="00:02:38.24"/><SPLIT distance="300" swimtime="00:04:01.11"/></SPLITS></RESULT><RESULT eventid="7" heatid="89" lane="5" points="387" resultid="669" swimtime="00:03:10.60"><SPLITS><SPLIT distance="50" swimtime="00:00:43.37"/><SPLIT distance="100" swimtime="00:01:32.91"/><SPLIT distance="150" swimtime="00:02:21.76"/></SPLITS></RESULT><RESULT eventid="9" heatid="120" lane="3" points="396" resultid="906" swimtime="00:00:32.23"><SPLITS/></RESULT><RESULT eventid="11" heatid="170" lane="8" points="401" resultid="1290" swimtime="00:02:50.92"><SPLITS><SPLIT distance="50" swimtime="00:00:38.32"/><SPLIT distance="100" swimtime="00:01:01.24"/><SPLIT distance="150" swimtime="00:02:13.43"/></SPLITS></RESULT><RESULT eventid="13" heatid="203" lane="2" points="331" resultid="1537" swimtime="00:01:23.04"><SPLITS><SPLIT distance="50" swimtime="00:00:40.24"/></SPLITS></RESULT><RESULT eventid="29" heatid="302" lane="8" points="395" resultid="2252" swimtime="00:02:33.94"><SPLITS><SPLIT distance="50" swimtime="00:00:34.74"/><SPLIT distance="100" swimtime="00:01:13.45"/><SPLIT distance="150" swimtime="00:01:55.59"/></SPLITS></RESULT><RESULT eventid="31" heatid="340" lane="2" points="375" resultid="2532" swimtime="00:01:28.88"><SPLITS><SPLIT distance="50" swimtime="00:00:42.01"/></SPLITS></RESULT><RESULT eventid="37" heatid="407" lane="3" points="376" resultid="3033" swimtime="00:02:50.84"><SPLITS><SPLIT distance="50" swimtime="00:00:40.67"/><SPLIT distance="100" swimtime="00:01:23.84"/><SPLIT distance="150" swimtime="00:02:08.53"/></SPLITS></RESULT><RESULT eventid="41" heatid="477" lane="1" points="420" resultid="3563" swimtime="00:05:55.54"><SPLITS><SPLIT distance="50" swimtime="00:00:37.96"/><SPLIT distance="100" swimtime="00:01:25.01"/><SPLIT distance="150" swimtime="00:02:12.01"/><SPLIT distance="200" swimtime="00:02:57.65"/><SPLIT distance="250" swimtime="00:03:46.91"/><SPLIT distance="300" swimtime="00:04:37.02"/><SPLIT distance="350" swimtime="00:05:16.73"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="360" birthdate="2011-01-01" firstname="Felizia" gender="F" lastname="Lemle" license="428886"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="50" lane="5" points="458" resultid="379" swimtime="00:05:06.64"><SPLITS><SPLIT distance="100" swimtime="00:01:12.33"/><SPLIT distance="200" swimtime="00:02:30.71"/><SPLIT distance="300" swimtime="00:03:49.88"/></SPLITS></RESULT><RESULT eventid="5" heatid="69" lane="8" points="361" resultid="519" swimtime="00:01:17.85"><SPLITS><SPLIT distance="50" swimtime="00:00:35.45"/></SPLITS></RESULT><RESULT eventid="11" heatid="172" lane="3" points="459" resultid="1301" swimtime="00:02:43.40"><SPLITS><SPLIT distance="50" swimtime="00:00:35.37"/><SPLIT distance="100" swimtime="00:01:16.28"/><SPLIT distance="150" swimtime="00:02:06.35"/></SPLITS></RESULT><RESULT eventid="13" heatid="207" lane="3" points="426" resultid="1570" swimtime="00:01:16.32"><SPLITS><SPLIT distance="50" swimtime="00:00:37.03"/></SPLITS></RESULT><RESULT eventid="27" heatid="271" lane="7" points="455" resultid="2016" swimtime="00:00:35.07"><SPLITS/></RESULT><RESULT eventid="29" heatid="304" lane="2" points="445" resultid="2262" swimtime="00:02:27.96"><SPLITS><SPLIT distance="50" swimtime="00:00:33.38"/><SPLIT distance="100" swimtime="00:01:10.79"/><SPLIT distance="150" swimtime="00:01:49.85"/></SPLITS></RESULT><RESULT eventid="35" heatid="380" lane="8" points="394" resultid="2835" swimtime="00:00:33.30"><SPLITS/></RESULT><RESULT eventid="37" heatid="410" lane="5" points="438" resultid="3059" swimtime="00:02:42.32"><SPLITS><SPLIT distance="50" swimtime="00:00:36.92"/><SPLIT distance="100" swimtime="00:01:17.86"/><SPLIT distance="150" swimtime="00:02:00.71"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="365" birthdate="2009-01-01" firstname="Antonia" gender="F" lastname="Hölzer" license="418054"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="51" lane="2" points="503" resultid="384" swimtime="00:04:57.06"><SPLITS><SPLIT distance="100" swimtime="00:01:10.00"/><SPLIT distance="200" swimtime="00:02:26.18"/><SPLIT distance="300" swimtime="00:03:43.14"/></SPLITS></RESULT><RESULT eventid="5" heatid="67" lane="5" points="332" resultid="500" swimtime="00:01:20.10"><SPLITS><SPLIT distance="50" swimtime="00:00:36.33"/></SPLITS></RESULT><RESULT eventid="11" heatid="172" lane="2" points="468" resultid="1300" swimtime="00:02:42.39"><SPLITS><SPLIT distance="50" swimtime="00:00:36.85"/><SPLIT distance="100" swimtime="00:01:14.58"/><SPLIT distance="150" swimtime="00:02:06.53"/></SPLITS></RESULT><RESULT eventid="13" heatid="208" lane="5" points="535" resultid="1579" swimtime="00:01:10.73"><SPLITS><SPLIT distance="50" swimtime="00:00:35.11"/></SPLITS></RESULT><RESULT eventid="27" heatid="272" lane="8" points="479" resultid="2024" swimtime="00:00:34.48"><SPLITS/></RESULT><RESULT eventid="29" heatid="304" lane="4" points="503" resultid="2264" swimtime="00:02:22.01"><SPLITS><SPLIT distance="50" swimtime="00:00:32.22"/><SPLIT distance="100" swimtime="00:01:08.84"/><SPLIT distance="150" swimtime="00:01:45.34"/></SPLITS></RESULT><RESULT eventid="37" heatid="412" lane="6" points="545" resultid="3076" swimtime="00:02:30.97"><SPLITS><SPLIT distance="100" swimtime="00:01:13.35"/></SPLITS></RESULT><RESULT eventid="39" heatid="446" lane="8" points="451" resultid="3335" swimtime="00:01:07.39"><SPLITS><SPLIT distance="50" swimtime="00:00:33.01"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="371" birthdate="2009-01-01" firstname="Ida" gender="F" lastname="Pfeuffer" license="407068"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="52" lane="1" points="497" resultid="390" swimtime="00:04:58.41"><SPLITS><SPLIT distance="100" swimtime="00:01:08.37"/><SPLIT distance="200" swimtime="00:02:24.62"/><SPLIT distance="300" swimtime="00:03:42.22"/></SPLITS></RESULT><RESULT eventid="5" heatid="69" lane="3" points="418" resultid="514" swimtime="00:01:14.16"><SPLITS><SPLIT distance="50" swimtime="00:00:34.80"/></SPLITS></RESULT><RESULT eventid="9" heatid="129" lane="6" points="513" resultid="980" swimtime="00:00:29.56"><SPLITS/></RESULT><RESULT eventid="15" heatid="227" lane="1" points="506" resultid="1716" swimtime="00:19:15.02"><SPLITS><SPLIT distance="100" swimtime="00:01:09.90"/><SPLIT distance="200" swimtime="00:02:25.02"/><SPLIT distance="300" swimtime="00:03:40.31"/><SPLIT distance="400" swimtime="00:04:56.99"/><SPLIT distance="500" swimtime="00:06:14.63"/><SPLIT distance="600" swimtime="00:07:32.40"/><SPLIT distance="700" swimtime="00:08:50.73"/><SPLIT distance="800" swimtime="00:10:09.89"/><SPLIT distance="900" swimtime="00:11:28.22"/><SPLIT distance="1000" swimtime="00:12:46.62"/><SPLIT distance="1100" swimtime="00:14:05.07"/><SPLIT distance="1200" swimtime="00:15:24.04"/><SPLIT distance="1300" swimtime="00:16:42.95"/><SPLIT distance="1400" swimtime="00:18:00.54"/></SPLITS></RESULT><RESULT eventid="29" heatid="306" lane="4" points="536" resultid="2278" swimtime="00:02:19.00"><SPLITS><SPLIT distance="50" swimtime="00:00:31.90"/><SPLIT distance="100" swimtime="00:01:06.83"/><SPLIT distance="150" swimtime="00:01:43.57"/></SPLITS></RESULT><RESULT eventid="33" heatid="359" lane="4" points="383" resultid="2670" swimtime="00:02:47.67"><SPLITS><SPLIT distance="50" swimtime="00:00:33.74"/><SPLIT distance="100" swimtime="00:01:15.61"/><SPLIT distance="150" swimtime="00:02:01.38"/></SPLITS></RESULT><RESULT eventid="35" heatid="379" lane="5" points="414" resultid="2824" swimtime="00:00:32.76"><SPLITS/></RESULT><RESULT eventid="39" heatid="449" lane="8" points="528" resultid="3357" swimtime="00:01:03.97"><SPLITS><SPLIT distance="50" swimtime="00:00:31.01"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="373" birthdate="2007-01-01" firstname="Sina" gender="F" lastname="Friedrich" license="439667"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="52" lane="3" points="597" resultid="392" swimtime="00:04:40.67"><SPLITS><SPLIT distance="100" swimtime="00:01:07.89"/><SPLIT distance="200" swimtime="00:02:17.71"/><SPLIT distance="300" swimtime="00:03:29.59"/></SPLITS></RESULT><RESULT eventid="9" heatid="130" lane="3" points="555" resultid="985" swimtime="00:00:28.79"><SPLITS/></RESULT><RESULT eventid="11" heatid="171" lane="4" points="505" resultid="1294" swimtime="00:02:38.35"><SPLITS><SPLIT distance="50" swimtime="00:00:34.19"/><SPLIT distance="100" swimtime="00:01:16.83"/><SPLIT distance="150" swimtime="00:02:05.14"/></SPLITS></RESULT><RESULT eventid="15" heatid="227" lane="7" points="552" resultid="1722" swimtime="00:18:41.57"><SPLITS><SPLIT distance="100" swimtime="00:01:11.83"/><SPLIT distance="200" swimtime="00:02:27.39"/><SPLIT distance="300" swimtime="00:03:42.72"/><SPLIT distance="400" swimtime="00:04:57.81"/><SPLIT distance="500" swimtime="00:06:12.72"/><SPLIT distance="600" swimtime="00:07:28.29"/><SPLIT distance="700" swimtime="00:08:43.35"/><SPLIT distance="800" swimtime="00:09:58.34"/><SPLIT distance="900" swimtime="00:11:13.05"/><SPLIT distance="1000" swimtime="00:12:28.06"/><SPLIT distance="1100" swimtime="00:13:43.31"/><SPLIT distance="1200" swimtime="00:14:59.30"/><SPLIT distance="1300" swimtime="00:16:14.74"/><SPLIT distance="1400" swimtime="00:17:29.80"/></SPLITS></RESULT><RESULT eventid="29" heatid="307" lane="6" points="633" resultid="2288" swimtime="00:02:11.58"><SPLITS><SPLIT distance="50" swimtime="00:00:30.93"/><SPLIT distance="100" swimtime="00:01:04.33"/><SPLIT distance="150" swimtime="00:01:38.53"/></SPLITS></RESULT><RESULT eventid="35" heatid="379" lane="3" points="396" resultid="2822" swimtime="00:00:33.26"><SPLITS/></RESULT><RESULT eventid="39" heatid="450" lane="6" points="589" resultid="3363" swimtime="00:01:01.68"><SPLITS><SPLIT distance="50" swimtime="00:00:29.96"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="374" birthdate="2010-01-01" firstname="Elisabeth" gender="F" lastname="Strecker" license="406754"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="52" lane="4" points="592" resultid="393" swimtime="00:04:41.54"><SPLITS><SPLIT distance="100" swimtime="00:01:06.81"/><SPLIT distance="200" swimtime="00:02:18.31"/><SPLIT distance="300" swimtime="00:03:30.55"/></SPLITS></RESULT><RESULT eventid="5" heatid="70" lane="5" points="477" resultid="524" swimtime="00:01:11.00"><SPLITS><SPLIT distance="50" swimtime="00:00:33.00"/></SPLITS></RESULT><RESULT eventid="9" heatid="131" lane="2" points="565" resultid="991" swimtime="00:00:28.62"><SPLITS/></RESULT><RESULT eventid="11" heatid="174" lane="8" points="527" resultid="1322" swimtime="00:02:36.07"><SPLITS><SPLIT distance="50" swimtime="00:00:33.62"/><SPLIT distance="100" swimtime="00:01:13.08"/><SPLIT distance="150" swimtime="00:02:02.37"/></SPLITS></RESULT><RESULT eventid="15" heatid="227" lane="3" points="536" resultid="1718" swimtime="00:18:52.83"><SPLITS><SPLIT distance="100" swimtime="00:01:09.00"/><SPLIT distance="200" swimtime="00:02:23.28"/><SPLIT distance="300" swimtime="00:03:38.00"/><SPLIT distance="400" swimtime="00:04:53.61"/><SPLIT distance="500" swimtime="00:06:09.21"/><SPLIT distance="600" swimtime="00:07:24.83"/><SPLIT distance="700" swimtime="00:08:40.88"/><SPLIT distance="800" swimtime="00:09:57.13"/><SPLIT distance="900" swimtime="00:11:13.24"/><SPLIT distance="1000" swimtime="00:12:29.92"/><SPLIT distance="1100" swimtime="00:13:47.15"/><SPLIT distance="1200" swimtime="00:15:04.57"/><SPLIT distance="1300" swimtime="00:16:21.70"/><SPLIT distance="1400" swimtime="00:17:37.95"/></SPLITS></RESULT><RESULT eventid="29" heatid="307" lane="5" points="612" resultid="2287" swimtime="00:02:13.04"><SPLITS><SPLIT distance="50" swimtime="00:00:30.97"/><SPLIT distance="100" swimtime="00:01:04.42"/><SPLIT distance="150" swimtime="00:01:39.00"/></SPLITS></RESULT><RESULT eventid="39" heatid="450" lane="5" points="588" resultid="3362" swimtime="00:01:01.69"><SPLITS><SPLIT distance="50" swimtime="00:00:29.89"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="375" birthdate="2008-01-01" firstname="Anouk" gender="F" lastname="Walther" license="346945"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="52" lane="5" points="605" resultid="394" swimtime="00:04:39.48"><SPLITS><SPLIT distance="100" swimtime="00:01:06.27"/><SPLIT distance="200" swimtime="00:02:17.35"/><SPLIT distance="300" swimtime="00:03:28.84"/></SPLITS></RESULT><RESULT eventid="5" heatid="71" lane="8" points="464" resultid="535" swimtime="00:01:11.64"><SPLITS><SPLIT distance="50" swimtime="00:00:33.72"/></SPLITS></RESULT><RESULT eventid="11" heatid="173" lane="4" points="587" resultid="1310" swimtime="00:02:30.58"><SPLITS><SPLIT distance="50" swimtime="00:00:31.38"/><SPLIT distance="100" swimtime="00:01:11.26"/><SPLIT distance="150" swimtime="00:01:57.51"/></SPLITS></RESULT><RESULT eventid="15" heatid="227" lane="4" points="631" resultid="1719" swimtime="00:17:52.98"><SPLITS><SPLIT distance="100" swimtime="00:01:07.20"/><SPLIT distance="200" swimtime="00:02:19.57"/><SPLIT distance="300" swimtime="00:03:31.66"/><SPLIT distance="400" swimtime="00:04:43.85"/><SPLIT distance="500" swimtime="00:05:55.95"/><SPLIT distance="600" swimtime="00:07:06.77"/><SPLIT distance="700" swimtime="00:08:18.57"/><SPLIT distance="800" swimtime="00:09:29.91"/><SPLIT distance="900" swimtime="00:10:41.89"/><SPLIT distance="1000" swimtime="00:11:53.93"/><SPLIT distance="1100" swimtime="00:13:06.05"/><SPLIT distance="1200" swimtime="00:14:18.53"/><SPLIT distance="1300" swimtime="00:15:30.23"/><SPLIT distance="1400" swimtime="00:16:42.17"/></SPLITS></RESULT><RESULT eventid="29" heatid="307" lane="2" points="554" resultid="2284" swimtime="00:02:17.51"><SPLITS><SPLIT distance="50" swimtime="00:00:31.63"/><SPLIT distance="100" swimtime="00:01:06.61"/><SPLIT distance="150" swimtime="00:01:42.25"/></SPLITS></RESULT><RESULT eventid="33" heatid="360" lane="6" points="515" resultid="2680" swimtime="00:02:31.92"><SPLITS><SPLIT distance="50" swimtime="00:00:32.67"/><SPLIT distance="100" swimtime="00:01:10.72"/><SPLIT distance="150" swimtime="00:01:50.78"/></SPLITS></RESULT><RESULT eventid="41" heatid="478" lane="3" points="588" resultid="3572" swimtime="00:05:17.93"><SPLITS><SPLIT distance="50" swimtime="00:00:32.64"/><SPLIT distance="100" swimtime="00:01:09.98"/><SPLIT distance="150" swimtime="00:01:52.08"/><SPLIT distance="200" swimtime="00:02:32.66"/><SPLIT distance="250" swimtime="00:03:19.73"/><SPLIT distance="300" swimtime="00:04:06.69"/><SPLIT distance="350" swimtime="00:04:43.21"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="378" birthdate="2011-01-01" firstname="Michelle" gender="F" lastname="Möbus" license="423840"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="52" lane="8" points="501" resultid="397" swimtime="00:04:57.55"><SPLITS><SPLIT distance="100" swimtime="00:01:09.87"/><SPLIT distance="200" swimtime="00:02:25.34"/><SPLIT distance="300" swimtime="00:03:42.26"/></SPLITS></RESULT><RESULT eventid="5" heatid="71" lane="1" points="485" resultid="528" swimtime="00:01:10.58"><SPLITS><SPLIT distance="50" swimtime="00:00:33.09"/></SPLITS></RESULT><RESULT eventid="11" heatid="173" lane="8" points="484" resultid="1314" swimtime="00:02:40.57"><SPLITS><SPLIT distance="50" swimtime="00:00:33.59"/><SPLIT distance="100" swimtime="00:01:15.13"/><SPLIT distance="150" swimtime="00:02:05.14"/></SPLITS></RESULT><RESULT eventid="13" heatid="208" lane="8" points="443" resultid="1582" swimtime="00:01:15.36"><SPLITS><SPLIT distance="50" swimtime="00:00:37.18"/></SPLITS></RESULT><RESULT eventid="29" heatid="306" lane="2" points="517" resultid="2276" swimtime="00:02:20.69"><SPLITS><SPLIT distance="50" swimtime="00:00:32.32"/><SPLIT distance="100" swimtime="00:01:07.52"/><SPLIT distance="150" swimtime="00:01:44.47"/></SPLITS></RESULT><RESULT eventid="33" heatid="360" lane="2" points="413" resultid="2676" swimtime="00:02:43.50"><SPLITS><SPLIT distance="50" swimtime="00:00:34.33"/><SPLIT distance="100" swimtime="00:01:14.05"/><SPLIT distance="150" swimtime="00:01:59.60"/></SPLITS></RESULT><RESULT eventid="35" heatid="381" lane="2" points="433" resultid="2837" swimtime="00:00:32.27"><SPLITS/></RESULT><RESULT eventid="37" heatid="411" lane="3" points="466" resultid="3065" swimtime="00:02:39.09"><SPLITS><SPLIT distance="100" swimtime="00:01:17.73"/></SPLITS></RESULT><RESULT eventid="41" heatid="478" lane="1" points="482" resultid="3570" swimtime="00:05:39.51"><SPLITS><SPLIT distance="50" swimtime="00:00:34.61"/><SPLIT distance="100" swimtime="00:01:16.14"/><SPLIT distance="150" swimtime="00:02:00.32"/><SPLIT distance="200" swimtime="00:02:43.12"/><SPLIT distance="250" swimtime="00:03:34.72"/><SPLIT distance="300" swimtime="00:04:25.64"/><SPLIT distance="350" swimtime="00:05:03.57"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="392" birthdate="2014-01-01" firstname="Jinqian" gender="M" lastname="Zhuang" license="481423"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="55" lane="6" points="202" resultid="415" swimtime="00:06:14.87"><SPLITS><SPLIT distance="100" swimtime="00:01:29.76"/><SPLIT distance="200" swimtime="00:03:08.66"/><SPLIT distance="300" swimtime="00:04:44.84"/></SPLITS></RESULT><RESULT eventid="8" heatid="93" lane="3" points="173" resultid="699" swimtime="00:03:46.03"><SPLITS><SPLIT distance="50" swimtime="00:00:54.27"/><SPLIT distance="100" swimtime="00:01:51.91"/><SPLIT distance="150" swimtime="00:02:51.73"/></SPLITS></RESULT><RESULT eventid="12" heatid="177" lane="1" points="172" resultid="1336" swimtime="00:03:24.91"><SPLITS><SPLIT distance="50" swimtime="00:00:49.62"/><SPLIT distance="100" swimtime="00:02:48.36"/><SPLIT distance="150" swimtime="00:02:40.30"/></SPLITS></RESULT><RESULT eventid="14" heatid="216" lane="1" points="149" resultid="1635" swimtime="00:01:37.18"><SPLITS><SPLIT distance="50" swimtime="00:00:47.79"/></SPLITS></RESULT><RESULT eventid="28" heatid="278" lane="6" points="142" resultid="2066" swimtime="00:00:45.35"><SPLITS/></RESULT><RESULT eventid="30" heatid="312" lane="2" points="193" resultid="2320" swimtime="00:02:56.26"><SPLITS><SPLIT distance="50" swimtime="00:00:39.50"/><SPLIT distance="100" swimtime="00:01:24.94"/><SPLIT distance="150" swimtime="00:02:11.72"/></SPLITS></RESULT><RESULT eventid="36" heatid="384" lane="4" points="121" resultid="2858" swimtime="00:00:44.96"><SPLITS/></RESULT><RESULT eventid="40" heatid="457" lane="4" points="188" resultid="3416" swimtime="00:01:21.70"><SPLITS><SPLIT distance="50" swimtime="00:00:39.36"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="400" birthdate="2015-01-01" firstname="Lukas" gender="M" lastname="Wällisch" license="479246"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="57" lane="1" points="238" resultid="426" swimtime="00:05:54.94"><SPLITS><SPLIT distance="100" swimtime="00:01:24.56"/><SPLIT distance="200" swimtime="00:02:56.37"/><SPLIT distance="300" swimtime="00:04:27.12"/></SPLITS></RESULT><RESULT eventid="6" heatid="73" lane="1" points="140" resultid="544" swimtime="00:01:35.12"><SPLITS><SPLIT distance="50" swimtime="00:00:44.56"/></SPLITS></RESULT><RESULT eventid="12" heatid="178" lane="5" points="221" resultid="1346" swimtime="00:03:08.45"><SPLITS><SPLIT distance="50" swimtime="00:00:42.76"/><SPLIT distance="100" swimtime="00:01:31.98"/><SPLIT distance="150" swimtime="00:02:26.07"/></SPLITS></RESULT><RESULT eventid="14" heatid="218" lane="5" points="186" resultid="1655" swimtime="00:01:30.27"><SPLITS><SPLIT distance="50" swimtime="00:00:45.14"/></SPLITS></RESULT><RESULT eventid="32" heatid="349" lane="5" points="175" resultid="2601" swimtime="00:01:41.53"><SPLITS><SPLIT distance="50" swimtime="00:00:48.09"/></SPLITS></RESULT><RESULT eventid="36" heatid="388" lane="1" points="150" resultid="2886" swimtime="00:00:41.84"><SPLITS/></RESULT><RESULT eventid="40" heatid="461" lane="3" points="207" resultid="3446" swimtime="00:01:19.11"><SPLITS><SPLIT distance="50" swimtime="00:00:37.08"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="402" birthdate="2009-01-01" firstname="Eric" gender="M" lastname="Lahner" license="409141"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="57" lane="3" points="270" resultid="428" swimtime="00:05:40.34"><SPLITS><SPLIT distance="100" swimtime="00:01:17.72"/><SPLIT distance="200" swimtime="00:02:41.53"/><SPLIT distance="300" swimtime="00:04:12.68"/></SPLITS></RESULT><RESULT eventid="10" heatid="147" lane="3" points="359" resultid="1108" swimtime="00:00:29.42"><SPLITS/></RESULT><RESULT eventid="14" heatid="221" lane="8" points="281" resultid="1681" swimtime="00:01:18.76"><SPLITS><SPLIT distance="50" swimtime="00:00:37.94"/></SPLITS></RESULT><RESULT eventid="28" heatid="283" lane="4" points="259" resultid="2104" swimtime="00:00:37.18"><SPLITS/></RESULT><RESULT eventid="30" heatid="318" lane="6" points="298" resultid="2371" swimtime="00:02:32.66"><SPLITS><SPLIT distance="50" swimtime="00:00:32.54"/><SPLIT distance="100" swimtime="00:01:11.46"/><SPLIT distance="150" swimtime="00:01:53.53"/></SPLITS></RESULT><RESULT eventid="36" heatid="393" lane="2" points="333" resultid="2927" swimtime="00:00:32.12"><SPLITS/></RESULT><RESULT eventid="38" heatid="417" lane="1" points="272" resultid="3107" swimtime="00:02:52.64"><SPLITS><SPLIT distance="50" swimtime="00:00:38.87"/><SPLIT distance="100" swimtime="00:01:21.79"/><SPLIT distance="150" swimtime="00:02:08.97"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="414" birthdate="2012-01-01" firstname="Felix" gender="M" lastname="Metz" license="435209"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="59" lane="3" points="428" resultid="443" swimtime="00:04:51.98"><SPLITS><SPLIT distance="100" swimtime="00:01:09.13"/><SPLIT distance="200" swimtime="00:02:23.51"/><SPLIT distance="300" swimtime="00:03:38.48"/></SPLITS></RESULT><RESULT eventid="6" heatid="73" lane="4" points="277" resultid="547" swimtime="00:01:15.85"><SPLITS><SPLIT distance="50" swimtime="00:00:35.02"/></SPLITS></RESULT><RESULT eventid="10" heatid="150" lane="1" points="378" resultid="1130" swimtime="00:00:28.90"><SPLITS/></RESULT><RESULT eventid="14" heatid="222" lane="7" points="292" resultid="1688" swimtime="00:01:17.70"><SPLITS><SPLIT distance="50" swimtime="00:00:37.77"/></SPLITS></RESULT><RESULT eventid="16" heatid="229" lane="7" points="404" resultid="1731" swimtime="00:19:37.80"><SPLITS><SPLIT distance="100" swimtime="00:01:12.67"/><SPLIT distance="200" swimtime="00:02:30.76"/><SPLIT distance="300" swimtime="00:03:49.61"/><SPLIT distance="400" swimtime="00:05:09.06"/><SPLIT distance="500" swimtime="00:06:28.47"/><SPLIT distance="600" swimtime="00:07:47.63"/><SPLIT distance="700" swimtime="00:09:07.21"/><SPLIT distance="800" swimtime="00:10:26.15"/><SPLIT distance="900" swimtime="00:11:44.94"/><SPLIT distance="1000" swimtime="00:13:03.94"/><SPLIT distance="1100" swimtime="00:14:22.88"/><SPLIT distance="1200" swimtime="00:15:42.10"/><SPLIT distance="1300" swimtime="00:17:01.57"/><SPLIT distance="1400" swimtime="00:18:20.51"/></SPLITS></RESULT><RESULT eventid="30" heatid="322" lane="7" points="403" resultid="2402" swimtime="00:02:17.98"><SPLITS><SPLIT distance="50" swimtime="00:00:30.96"/><SPLIT distance="100" swimtime="00:01:06.56"/><SPLIT distance="150" swimtime="00:01:42.82"/></SPLITS></RESULT><RESULT eventid="36" heatid="392" lane="6" points="351" resultid="2923" swimtime="00:00:31.57"><SPLITS/></RESULT><RESULT eventid="40" heatid="469" lane="1" points="416" resultid="3506" swimtime="00:01:02.76"><SPLITS><SPLIT distance="50" swimtime="00:00:30.63"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="416" birthdate="2011-01-01" firstname="Kai" gender="M" lastname="Crazzolara" license="425766"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="59" lane="5" points="392" resultid="445" swimtime="00:05:00.47"><SPLITS><SPLIT distance="100" swimtime="00:01:11.83"/><SPLIT distance="200" swimtime="00:02:30.33"/><SPLIT distance="300" swimtime="00:03:48.05"/></SPLITS></RESULT><RESULT eventid="6" heatid="76" lane="5" points="311" resultid="571" swimtime="00:01:12.95"><SPLITS><SPLIT distance="50" swimtime="00:00:33.59"/></SPLITS></RESULT><RESULT eventid="10" heatid="149" lane="7" points="384" resultid="1128" swimtime="00:00:28.76"><SPLITS/></RESULT><RESULT eventid="12" heatid="186" lane="8" points="359" resultid="1411" swimtime="00:02:40.32"><SPLITS><SPLIT distance="50" swimtime="00:00:34.79"/><SPLIT distance="100" swimtime="00:01:16.87"/><SPLIT distance="150" swimtime="00:02:06.17"/></SPLITS></RESULT><RESULT eventid="16" heatid="229" lane="1" points="383" resultid="1726" swimtime="00:19:59.27"><SPLITS><SPLIT distance="100" swimtime="00:01:13.34"/><SPLIT distance="200" swimtime="00:02:34.68"/><SPLIT distance="300" swimtime="00:03:55.94"/><SPLIT distance="400" swimtime="00:05:17.82"/><SPLIT distance="500" swimtime="00:06:37.64"/><SPLIT distance="600" swimtime="00:07:57.81"/><SPLIT distance="700" swimtime="00:09:18.43"/><SPLIT distance="800" swimtime="00:10:38.99"/><SPLIT distance="900" swimtime="00:12:00.78"/><SPLIT distance="1000" swimtime="00:13:22.69"/><SPLIT distance="1100" swimtime="00:14:44.35"/><SPLIT distance="1200" swimtime="00:16:06.88"/><SPLIT distance="1300" swimtime="00:17:26.49"/><SPLIT distance="1400" swimtime="00:18:45.72"/></SPLITS></RESULT><RESULT eventid="28" heatid="283" lane="3" points="328" resultid="2103" swimtime="00:00:34.37"><SPLITS/></RESULT><RESULT eventid="30" heatid="321" lane="6" points="388" resultid="2393" swimtime="00:02:19.80"><SPLITS><SPLIT distance="50" swimtime="00:00:32.39"/><SPLIT distance="100" swimtime="00:01:09.12"/><SPLIT distance="150" swimtime="00:01:45.77"/></SPLITS></RESULT><RESULT eventid="40" heatid="468" lane="2" points="400" resultid="3499" swimtime="00:01:03.56"><SPLITS><SPLIT distance="50" swimtime="00:00:30.10"/></SPLITS></RESULT><RESULT eventid="42" heatid="479" lane="5" points="388" resultid="3581" swimtime="00:05:34.19"><SPLITS><SPLIT distance="50" swimtime="00:00:35.08"/><SPLIT distance="100" swimtime="00:01:16.75"/><SPLIT distance="150" swimtime="00:02:00.40"/><SPLIT distance="200" swimtime="00:02:43.22"/><SPLIT distance="250" swimtime="00:03:30.75"/><SPLIT distance="300" swimtime="00:04:19.56"/><SPLIT distance="350" swimtime="00:04:57.98"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="420" birthdate="2011-01-01" firstname="Michael" gender="M" lastname="Polubock" license="480832"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="60" lane="1" points="403" resultid="449" swimtime="00:04:57.72"><SPLITS><SPLIT distance="100" swimtime="00:01:11.31"/><SPLIT distance="200" swimtime="00:02:27.41"/><SPLIT distance="300" swimtime="00:03:43.34"/></SPLITS></RESULT><RESULT eventid="6" heatid="77" lane="8" points="332" resultid="582" swimtime="00:01:11.37"><SPLITS><SPLIT distance="50" swimtime="00:00:34.12"/></SPLITS></RESULT><RESULT eventid="10" heatid="149" lane="8" points="408" resultid="1129" swimtime="00:00:28.17"><SPLITS/></RESULT><RESULT eventid="12" heatid="186" lane="2" points="389" resultid="1405" swimtime="00:02:36.13"><SPLITS><SPLIT distance="50" swimtime="00:00:32.70"/><SPLIT distance="100" swimtime="00:01:14.35"/><SPLIT distance="150" swimtime="00:01:59.28"/></SPLITS></RESULT><RESULT eventid="30" heatid="321" lane="7" points="371" resultid="2394" swimtime="00:02:21.92"><SPLITS><SPLIT distance="50" swimtime="00:00:31.20"/><SPLIT distance="100" swimtime="00:01:07.72"/><SPLIT distance="150" swimtime="00:01:44.80"/></SPLITS></RESULT><RESULT eventid="32" heatid="352" lane="1" points="307" resultid="2620" swimtime="00:01:24.26"><SPLITS><SPLIT distance="50" swimtime="00:00:40.62"/></SPLITS></RESULT><RESULT eventid="36" heatid="394" lane="3" points="377" resultid="2936" swimtime="00:00:30.81"><SPLITS/></RESULT><RESULT eventid="40" heatid="469" lane="7" points="442" resultid="3512" swimtime="00:01:01.51"><SPLITS><SPLIT distance="50" swimtime="00:00:29.68"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="428" birthdate="1996-01-01" firstname="Alexander" gender="M" lastname="Klingert" license="169874"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="61" lane="2" points="459" resultid="457" swimtime="00:04:45.26"><SPLITS><SPLIT distance="100" swimtime="00:01:02.79"/><SPLIT distance="200" swimtime="00:02:14.97"/><SPLIT distance="300" swimtime="00:03:30.19"/></SPLITS></RESULT><RESULT eventid="12" heatid="189" lane="7" points="484" resultid="1433" swimtime="00:02:25.12"><SPLITS><SPLIT distance="50" swimtime="00:00:29.92"/><SPLIT distance="100" swimtime="00:01:08.10"/><SPLIT distance="150" swimtime="00:01:52.51"/></SPLITS></RESULT><RESULT eventid="14" heatid="225" lane="7" points="487" resultid="1710" swimtime="00:01:05.58"><SPLITS><SPLIT distance="50" swimtime="00:00:31.40"/></SPLITS></RESULT><RESULT eventid="30" heatid="324" lane="4" points="501" resultid="2414" swimtime="00:02:08.40"><SPLITS><SPLIT distance="50" swimtime="00:00:28.37"/><SPLIT distance="100" swimtime="00:00:59.79"/><SPLIT distance="150" swimtime="00:01:33.80"/></SPLITS></RESULT><RESULT eventid="40" heatid="475" lane="8" points="554" resultid="3559" swimtime="00:00:57.03"><SPLITS><SPLIT distance="50" swimtime="00:00:27.98"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="435" birthdate="2001-01-01" firstname="Philipp" gender="M" lastname="Harig" license="300003"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="62" lane="3" points="455" resultid="464" swimtime="00:04:46.00"><SPLITS><SPLIT distance="100" swimtime="00:01:03.22"/><SPLIT distance="200" swimtime="00:02:14.75"/><SPLIT distance="300" swimtime="00:03:29.90"/></SPLITS></RESULT><RESULT eventid="12" heatid="189" lane="2" points="464" resultid="1429" swimtime="00:02:27.20"><SPLITS><SPLIT distance="50" swimtime="00:00:30.81"/><SPLIT distance="100" swimtime="00:01:06.26"/><SPLIT distance="150" swimtime="00:01:52.93"/></SPLITS></RESULT><RESULT eventid="14" heatid="225" lane="1" points="460" resultid="1705" swimtime="00:01:06.84"><SPLITS><SPLIT distance="50" swimtime="00:00:31.71"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="463" birthdate="2004-01-01" firstname="Jana" gender="F" lastname="Birner" license="354619"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="5" heatid="71" lane="3" points="553" resultid="530" swimtime="00:01:07.59"><SPLITS><SPLIT distance="50" swimtime="00:00:31.43"/></SPLITS></RESULT><RESULT eventid="9" heatid="131" lane="1" points="554" resultid="990" swimtime="00:00:28.81"><SPLITS/></RESULT><RESULT eventid="35" heatid="382" lane="5" points="552" resultid="2848" swimtime="00:00:29.77"><SPLITS/></RESULT><RESULT eventid="39" heatid="450" lane="7" points="578" resultid="3364" swimtime="00:01:02.05"><SPLITS><SPLIT distance="50" swimtime="00:00:29.73"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="470" birthdate="2010-01-01" firstname="Paul" gender="M" lastname="Welker" license="416995"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="6" heatid="72" lane="6" points="192" resultid="541" swimtime="00:01:25.64"><SPLITS><SPLIT distance="50" swimtime="00:00:36.61"/></SPLITS></RESULT><RESULT eventid="10" heatid="148" lane="1" points="293" resultid="1114" swimtime="00:00:31.47"><SPLITS/></RESULT><RESULT eventid="12" heatid="181" lane="5" points="283" resultid="1370" swimtime="00:02:53.53"><SPLITS><SPLIT distance="50" swimtime="00:00:39.41"/><SPLIT distance="100" swimtime="00:01:26.25"/><SPLIT distance="150" swimtime="00:02:16.51"/></SPLITS></RESULT><RESULT eventid="30" heatid="320" lane="3" points="329" resultid="2384" swimtime="00:02:27.62"><SPLITS><SPLIT distance="50" swimtime="00:00:34.10"/><SPLIT distance="100" swimtime="00:01:11.46"/><SPLIT distance="150" swimtime="00:01:50.50"/></SPLITS></RESULT><RESULT eventid="32" heatid="352" lane="2" points="310" resultid="2621" swimtime="00:01:24.01"><SPLITS><SPLIT distance="50" swimtime="00:00:39.99"/></SPLITS></RESULT><RESULT eventid="36" heatid="392" lane="8" points="209" resultid="2925" swimtime="00:00:37.50"><SPLITS/></RESULT><RESULT eventid="40" heatid="467" lane="1" points="289" resultid="3491" swimtime="00:01:10.81"><SPLITS><SPLIT distance="50" swimtime="00:00:34.22"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="473" birthdate="2011-01-01" firstname="Samuel" gender="M" lastname="Jakubietz" license="436705"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="6" heatid="73" lane="3" points="189" resultid="546" swimtime="00:01:26.06"><SPLITS><SPLIT distance="50" swimtime="00:00:37.67"/></SPLITS></RESULT><RESULT eventid="10" heatid="146" lane="4" points="306" resultid="1101" swimtime="00:00:31.00"><SPLITS/></RESULT><RESULT eventid="12" heatid="182" lane="6" points="291" resultid="1379" swimtime="00:02:51.87"><SPLITS><SPLIT distance="50" swimtime="00:00:37.23"/><SPLIT distance="100" swimtime="00:01:23.28"/><SPLIT distance="150" swimtime="00:02:12.89"/></SPLITS></RESULT><RESULT eventid="28" heatid="282" lane="3" points="239" resultid="2095" swimtime="00:00:38.20"><SPLITS/></RESULT><RESULT eventid="30" heatid="322" lane="8" points="290" resultid="2403" swimtime="00:02:34.00"><SPLITS><SPLIT distance="50" swimtime="00:00:34.72"/><SPLIT distance="100" swimtime="00:01:13.50"/><SPLIT distance="150" swimtime="00:01:55.87"/></SPLITS></RESULT><RESULT eventid="36" heatid="391" lane="1" points="224" resultid="2910" swimtime="00:00:36.64"><SPLITS/></RESULT><RESULT eventid="40" heatid="466" lane="6" points="338" resultid="3488" swimtime="00:01:07.27"><SPLITS><SPLIT distance="50" swimtime="00:00:32.63"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="474" birthdate="2011-01-01" firstname="Eric" gender="M" lastname="Baumstark" license="444895"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="6" heatid="73" lane="6" points="205" resultid="548" swimtime="00:01:23.85"><SPLITS><SPLIT distance="50" swimtime="00:00:38.02"/></SPLITS></RESULT><RESULT eventid="10" heatid="145" lane="4" points="288" resultid="1093" swimtime="00:00:31.65"><SPLITS/></RESULT><RESULT eventid="12" heatid="179" lane="4" points="236" resultid="1353" swimtime="00:03:04.37"><SPLITS><SPLIT distance="50" swimtime="00:00:38.05"/><SPLIT distance="100" swimtime="00:01:25.61"/><SPLIT distance="150" swimtime="00:02:22.57"/></SPLITS></RESULT><RESULT eventid="28" heatid="280" lane="4" points="207" resultid="2080" swimtime="00:00:40.08"><SPLITS/></RESULT><RESULT eventid="30" heatid="318" lane="8" points="240" resultid="2373" swimtime="00:02:44.07"><SPLITS><SPLIT distance="50" swimtime="00:00:36.11"/><SPLIT distance="100" swimtime="00:01:18.09"/><SPLIT distance="150" swimtime="00:02:03.69"/></SPLITS></RESULT><RESULT eventid="36" heatid="391" lane="4" points="279" resultid="2913" swimtime="00:00:34.08"><SPLITS/></RESULT><RESULT eventid="40" heatid="465" lane="1" points="274" resultid="3475" swimtime="00:01:12.11"><SPLITS><SPLIT distance="50" swimtime="00:00:35.26"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="475" birthdate="2011-01-01" firstname="Henri" gender="M" lastname="Kiessig" license="447240"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="6" heatid="73" lane="7" points="161" resultid="549" swimtime="00:01:30.88"><SPLITS><SPLIT distance="50" swimtime="00:00:41.03"/></SPLITS></RESULT><RESULT eventid="10" heatid="144" lane="6" points="240" resultid="1087" swimtime="00:00:33.63"><SPLITS/></RESULT><RESULT eventid="14" heatid="218" lane="4" points="234" resultid="1654" swimtime="00:01:23.62"><SPLITS><SPLIT distance="50" swimtime="00:00:40.45"/></SPLITS></RESULT><RESULT eventid="28" heatid="283" lane="7" points="251" resultid="2107" swimtime="00:00:37.57"><SPLITS/></RESULT><RESULT eventid="30" heatid="316" lane="5" points="221" resultid="2354" swimtime="00:02:48.57"><SPLITS><SPLIT distance="50" swimtime="00:00:38.12"/><SPLIT distance="100" swimtime="00:01:21.10"/><SPLIT distance="150" swimtime="00:02:05.96"/></SPLITS></RESULT><RESULT eventid="36" heatid="390" lane="4" points="208" resultid="2905" swimtime="00:00:37.55"><SPLITS/></RESULT><RESULT eventid="40" heatid="464" lane="7" points="260" resultid="3473" swimtime="00:01:13.36"><SPLITS><SPLIT distance="50" swimtime="00:00:35.37"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="489" birthdate="2006-01-01" firstname="Richard" gender="M" lastname="Knecht" license="349713"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="6" heatid="77" lane="3" points="395" resultid="577" swimtime="00:01:07.35"><SPLITS><SPLIT distance="50" swimtime="00:00:31.51"/></SPLITS></RESULT><RESULT eventid="10" heatid="151" lane="7" points="424" resultid="1144" swimtime="00:00:27.83"><SPLITS/></RESULT><RESULT eventid="12" heatid="187" lane="6" points="389" resultid="1417" swimtime="00:02:36.14"><SPLITS><SPLIT distance="50" swimtime="00:00:31.33"/><SPLIT distance="100" swimtime="00:01:13.46"/><SPLIT distance="150" swimtime="00:02:01.38"/></SPLITS></RESULT><RESULT eventid="40" heatid="470" lane="8" resultid="3521" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="490" birthdate="1999-01-01" firstname="Jindrich" gender="M" lastname="Sedlacek" license="267952"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="6" heatid="77" lane="4" points="314" resultid="578" swimtime="00:01:12.69"><SPLITS><SPLIT distance="50" swimtime="00:00:34.23"/></SPLITS></RESULT><RESULT eventid="10" heatid="150" lane="7" points="383" resultid="1136" swimtime="00:00:28.79"><SPLITS/></RESULT><RESULT eventid="36" heatid="396" lane="6" points="357" resultid="2955" swimtime="00:00:31.37"><SPLITS/></RESULT><RESULT eventid="40" heatid="469" lane="6" points="417" resultid="3511" swimtime="00:01:02.68"><SPLITS><SPLIT distance="50" swimtime="00:00:29.73"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="497" birthdate="1997-01-01" firstname="Roland" gender="M" lastname="Hoffmann" license="237457"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="6" heatid="79" lane="1" points="489" resultid="590" swimtime="00:01:02.76"><SPLITS><SPLIT distance="50" swimtime="00:00:29.11"/></SPLITS></RESULT><RESULT eventid="10" heatid="156" lane="1" points="501" resultid="1176" swimtime="00:00:26.31"><SPLITS/></RESULT><RESULT eventid="30" heatid="324" lane="7" points="503" resultid="2417" swimtime="00:02:08.20"><SPLITS><SPLIT distance="50" swimtime="00:00:28.94"/><SPLIT distance="100" swimtime="00:01:00.98"/><SPLIT distance="150" swimtime="00:01:34.32"/></SPLITS></RESULT><RESULT eventid="36" heatid="399" lane="4" points="542" resultid="2977" swimtime="00:00:27.31"><SPLITS/></RESULT><RESULT eventid="40" heatid="475" lane="1" points="544" resultid="3552" swimtime="00:00:57.37"><SPLITS><SPLIT distance="50" swimtime="00:00:27.24"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="500" birthdate="2006-01-01" firstname="Paul" gender="M" lastname="Ziemainz" license="403946"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="6" heatid="80" lane="3" points="513" resultid="599" swimtime="00:01:01.74"><SPLITS><SPLIT distance="50" swimtime="00:00:28.61"/></SPLITS></RESULT><RESULT eventid="10" heatid="156" lane="3" points="509" resultid="1178" swimtime="00:00:26.18"><SPLITS/></RESULT><RESULT eventid="14" heatid="225" lane="6" points="480" resultid="1709" swimtime="00:01:05.86"><SPLITS><SPLIT distance="50" swimtime="00:00:31.46"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="516" birthdate="2007-01-01" firstname="Yasmin" gender="F" lastname="Yaser Salih" license="404986"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="9" heatid="113" lane="4" points="221" resultid="852" swimtime="00:00:39.12"><SPLITS/></RESULT><RESULT eventid="29" heatid="293" lane="7" points="195" resultid="2180" swimtime="00:03:14.57"><SPLITS><SPLIT distance="50" swimtime="00:00:42.63"/><SPLIT distance="100" swimtime="00:01:31.45"/><SPLIT distance="150" swimtime="00:02:24.29"/></SPLITS></RESULT><RESULT eventid="35" heatid="366" lane="2" points="129" resultid="2720" swimtime="00:00:48.23"><SPLITS/></RESULT><RESULT eventid="39" heatid="430" lane="6" points="199" resultid="3207" swimtime="00:01:28.53"><SPLITS><SPLIT distance="50" swimtime="00:00:41.80"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="517" birthdate="2010-01-01" firstname="Mia" gender="F" lastname="Schenk" license="436830"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="9" heatid="118" lane="5" points="364" resultid="892" swimtime="00:00:33.15"><SPLITS/></RESULT><RESULT eventid="11" heatid="165" lane="7" points="312" resultid="1249" swimtime="00:03:05.77"><SPLITS><SPLIT distance="50" swimtime="00:00:39.34"/><SPLIT distance="100" swimtime="00:01:30.24"/><SPLIT distance="150" swimtime="00:02:25.41"/></SPLITS></RESULT><RESULT eventid="13" heatid="202" lane="8" points="281" resultid="1535" swimtime="00:01:27.66"><SPLITS><SPLIT distance="50" swimtime="00:00:43.90"/></SPLITS></RESULT><RESULT eventid="27" heatid="266" lane="7" points="348" resultid="1978" swimtime="00:00:38.34"><SPLITS/></RESULT><RESULT eventid="29" heatid="298" lane="5" points="336" resultid="2218" swimtime="00:02:42.38"><SPLITS><SPLIT distance="50" swimtime="00:00:37.94"/><SPLIT distance="100" swimtime="00:01:20.56"/></SPLITS></RESULT><RESULT eventid="37" heatid="405" lane="4" points="280" resultid="3018" swimtime="00:03:08.39"><SPLITS><SPLIT distance="50" swimtime="00:00:44.79"/><SPLIT distance="100" swimtime="00:01:34.97"/><SPLIT distance="150" swimtime="00:02:23.66"/></SPLITS></RESULT><RESULT eventid="39" heatid="437" lane="8" points="328" resultid="3265" swimtime="00:01:14.97"><SPLITS><SPLIT distance="50" swimtime="00:00:36.56"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="518" birthdate="2009-01-01" firstname="Lina Malu" gender="F" lastname="Weßendorf" license="470858"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="9" heatid="118" lane="8" points="303" resultid="895" swimtime="00:00:35.22"><SPLITS/></RESULT><RESULT eventid="13" heatid="200" lane="7" points="221" resultid="1518" swimtime="00:01:34.88"><SPLITS><SPLIT distance="50" swimtime="00:00:46.63"/></SPLITS></RESULT><RESULT eventid="27" heatid="264" lane="1" points="246" resultid="1956" swimtime="00:00:43.03"><SPLITS/></RESULT><RESULT eventid="29" heatid="296" lane="8" points="278" resultid="2205" swimtime="00:02:53.00"><SPLITS><SPLIT distance="50" swimtime="00:00:38.62"/><SPLIT distance="100" swimtime="00:01:21.53"/><SPLIT distance="150" swimtime="00:02:08.30"/></SPLITS></RESULT><RESULT eventid="37" heatid="404" lane="2" points="250" resultid="3008" swimtime="00:03:15.69"><SPLITS><SPLIT distance="50" swimtime="00:00:46.00"/><SPLIT distance="100" swimtime="00:01:35.38"/><SPLIT distance="150" swimtime="00:02:26.34"/></SPLITS></RESULT><RESULT eventid="39" heatid="436" lane="2" points="299" resultid="3251" swimtime="00:01:17.29"><SPLITS><SPLIT distance="50" swimtime="00:00:36.59"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="519" birthdate="2012-01-01" firstname="Mathea" gender="F" lastname="Zentner" license="446975"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="9" heatid="119" lane="4" points="413" resultid="899" swimtime="00:00:31.78"><SPLITS/></RESULT><RESULT eventid="11" heatid="163" lane="1" points="298" resultid="1227" swimtime="00:03:08.78"><SPLITS><SPLIT distance="50" swimtime="00:00:39.94"/><SPLIT distance="100" swimtime="00:01:25.42"/><SPLIT distance="150" swimtime="00:02:27.20"/></SPLITS></RESULT><RESULT eventid="13" heatid="200" lane="6" resultid="1517" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="520" birthdate="2009-01-01" firstname="Elisabeth" gender="F" lastname="Lorenz" license="430176"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="9" heatid="119" lane="7" points="356" resultid="902" swimtime="00:00:33.39"><SPLITS/></RESULT><RESULT eventid="11" heatid="164" lane="5" points="280" resultid="1239" swimtime="00:03:12.77"><SPLITS><SPLIT distance="50" swimtime="00:00:40.32"/><SPLIT distance="100" swimtime="00:01:32.33"/><SPLIT distance="150" swimtime="00:02:27.62"/></SPLITS></RESULT><RESULT eventid="27" heatid="262" lane="4" points="268" resultid="1943" swimtime="00:00:41.81"><SPLITS/></RESULT><RESULT eventid="29" heatid="297" lane="3" points="299" resultid="2208" swimtime="00:02:48.84"><SPLITS><SPLIT distance="50" swimtime="00:00:38.72"/><SPLIT distance="100" swimtime="00:01:21.20"/><SPLIT distance="150" swimtime="00:02:06.99"/></SPLITS></RESULT><RESULT eventid="35" heatid="373" lane="8" points="256" resultid="2782" swimtime="00:00:38.46"><SPLITS/></RESULT><RESULT eventid="39" heatid="437" lane="3" points="323" resultid="3260" swimtime="00:01:15.33"><SPLITS><SPLIT distance="50" swimtime="00:00:35.83"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="521" birthdate="2007-01-01" firstname="Alba" gender="F" lastname="Warter Rubio" license="373291"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="9" heatid="120" lane="6" points="356" resultid="909" swimtime="00:00:33.37"><SPLITS/></RESULT><RESULT eventid="29" heatid="299" lane="5" points="304" resultid="2226" swimtime="00:02:47.87"><SPLITS><SPLIT distance="50" swimtime="00:00:36.20"/><SPLIT distance="100" swimtime="00:01:18.05"/><SPLIT distance="150" swimtime="00:02:03.45"/></SPLITS></RESULT><RESULT eventid="39" heatid="438" lane="4" points="337" resultid="3269" swimtime="00:01:14.29"><SPLITS><SPLIT distance="50" swimtime="00:00:34.27"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="526" birthdate="2010-01-01" firstname="Annika" gender="F" lastname="Zimmermann" license="416996"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="9" heatid="123" lane="6" resultid="933" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="13" heatid="203" lane="7" resultid="1542" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="27" heatid="267" lane="5" resultid="1984" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="29" heatid="299" lane="1" resultid="2222" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="37" heatid="407" lane="2" resultid="3032" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="39" heatid="438" lane="6" resultid="3271" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="530" birthdate="1999-01-01" firstname="Anna" gender="F" lastname="Pfretzschner" license="268769"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="9" heatid="128" lane="6" points="501" resultid="972" swimtime="00:00:29.80"><SPLITS/></RESULT><RESULT eventid="11" heatid="167" lane="1" points="354" resultid="1259" swimtime="00:02:58.17"><SPLITS><SPLIT distance="50" swimtime="00:00:35.45"/><SPLIT distance="100" swimtime="00:01:20.46"/><SPLIT distance="150" swimtime="00:02:15.83"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="534" birthdate="2008-01-01" firstname="Carla" gender="F" lastname="Primorac" license="392227"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="9" heatid="131" lane="7" points="599" resultid="995" swimtime="00:00:28.07"><SPLITS/></RESULT><RESULT eventid="11" heatid="173" lane="3" points="508" resultid="1309" swimtime="00:02:37.99"><SPLITS><SPLIT distance="50" swimtime="00:00:34.36"/><SPLIT distance="100" swimtime="00:01:15.22"/><SPLIT distance="150" swimtime="00:02:02.94"/></SPLITS></RESULT><RESULT eventid="29" heatid="307" lane="8" points="534" resultid="2290" swimtime="00:02:19.23"><SPLITS><SPLIT distance="50" swimtime="00:00:31.85"/><SPLIT distance="100" swimtime="00:01:06.59"/><SPLIT distance="150" swimtime="00:01:42.90"/></SPLITS></RESULT><RESULT eventid="35" heatid="381" lane="4" points="406" resultid="2839" swimtime="00:00:32.98"><SPLITS/></RESULT><RESULT eventid="39" heatid="450" lane="1" points="570" resultid="3358" swimtime="00:01:02.35"><SPLITS><SPLIT distance="50" swimtime="00:00:29.98"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="542" birthdate="2011-01-01" firstname="Finn" gender="M" lastname="Fritzsch" license="460136"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="10" heatid="138" lane="5" points="161" resultid="1041" swimtime="00:00:38.42"><SPLITS/></RESULT><RESULT eventid="14" heatid="213" lane="7" points="122" resultid="1619" swimtime="00:01:44.03"><SPLITS><SPLIT distance="50" swimtime="00:00:51.17"/></SPLITS></RESULT><RESULT eventid="28" heatid="275" lane="7" points="118" resultid="2045" swimtime="00:00:48.29"><SPLITS/></RESULT><RESULT eventid="30" heatid="312" lane="6" points="147" resultid="2324" swimtime="00:03:13.14"><SPLITS><SPLIT distance="50" swimtime="00:00:42.97"/><SPLIT distance="100" swimtime="00:01:30.26"/><SPLIT distance="150" swimtime="00:02:23.08"/></SPLITS></RESULT><RESULT eventid="40" heatid="457" lane="7" points="137" resultid="3419" swimtime="00:01:30.82"><SPLITS><SPLIT distance="50" swimtime="00:00:41.47"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="543" birthdate="2014-01-01" firstname="Timo" gender="M" lastname="Stecher" license="462915"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="10" heatid="139" lane="2" points="164" resultid="1045" swimtime="00:00:38.17"><SPLITS/></RESULT><RESULT comment="16:06 Der Sportler hat die Teilstrecke Rücken nicht in Rückenlage beendet" eventid="12" heatid="176" lane="1" resultid="1328" status="DSQ" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="14" heatid="213" lane="5" points="120" resultid="1617" swimtime="00:01:44.33"><SPLITS><SPLIT distance="50" swimtime="00:00:51.52"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="544" birthdate="2012-01-01" firstname="Oskar" gender="M" lastname="Kiessig" license="460137"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="10" heatid="139" lane="8" points="151" resultid="1051" swimtime="00:00:39.24"><SPLITS/></RESULT><RESULT eventid="14" heatid="212" lane="5" points="104" resultid="1609" swimtime="00:01:49.59"><SPLITS><SPLIT distance="50" swimtime="00:00:53.98"/></SPLITS></RESULT><RESULT eventid="28" heatid="277" lane="1" points="109" resultid="2054" swimtime="00:00:49.62"><SPLITS/></RESULT><RESULT eventid="40" heatid="456" lane="5" points="145" resultid="3410" swimtime="00:01:29.11"><SPLITS><SPLIT distance="50" swimtime="00:00:43.67"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="549" birthdate="2011-01-01" firstname="Dennes" gender="M" lastname="Ying" license="446974"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="10" heatid="146" lane="1" points="300" resultid="1098" swimtime="00:00:31.23"><SPLITS/></RESULT><RESULT eventid="12" heatid="180" lane="1" points="217" resultid="1358" swimtime="00:03:09.70"><SPLITS><SPLIT distance="50" swimtime="00:00:39.23"/><SPLIT distance="100" swimtime="00:01:28.22"/><SPLIT distance="150" swimtime="00:02:24.79"/></SPLITS></RESULT><RESULT eventid="28" heatid="280" lane="5" points="254" resultid="2081" swimtime="00:00:37.40"><SPLITS/></RESULT><RESULT eventid="32" heatid="351" lane="7" points="240" resultid="2618" swimtime="00:01:31.47"><SPLITS><SPLIT distance="50" swimtime="00:00:41.74"/></SPLITS></RESULT><RESULT eventid="36" heatid="390" lane="1" points="184" resultid="2902" swimtime="00:00:39.10"><SPLITS/></RESULT><RESULT eventid="40" heatid="464" lane="8" points="252" resultid="3474" swimtime="00:01:14.17"><SPLITS><SPLIT distance="50" swimtime="00:00:34.58"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="550" birthdate="2010-01-01" firstname="Ruben" gender="M" lastname="Riehle Mendez" license="423317"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="10" heatid="146" lane="7" points="299" resultid="1104" swimtime="00:00:31.27"><SPLITS/></RESULT><RESULT eventid="14" heatid="220" lane="2" points="210" resultid="1668" swimtime="00:01:26.76"><SPLITS><SPLIT distance="50" swimtime="00:00:41.36"/></SPLITS></RESULT><RESULT comment="09:41 Start vor dem Startsignal" eventid="28" heatid="280" lane="6" resultid="2082" status="DSQ" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="30" heatid="315" lane="6" points="195" resultid="2347" swimtime="00:02:55.61"><SPLITS><SPLIT distance="50" swimtime="00:00:38.54"/><SPLIT distance="100" swimtime="00:01:22.28"/><SPLIT distance="150" swimtime="00:02:09.61"/></SPLITS></RESULT><RESULT eventid="38" heatid="416" lane="6" points="216" resultid="3104" swimtime="00:03:06.50"><SPLITS><SPLIT distance="50" swimtime="00:00:41.71"/><SPLIT distance="100" swimtime="00:01:28.67"/><SPLIT distance="150" swimtime="00:02:18.49"/></SPLITS></RESULT><RESULT eventid="40" heatid="464" lane="2" points="210" resultid="3468" swimtime="00:01:18.80"><SPLITS><SPLIT distance="50" swimtime="00:00:36.34"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="551" birthdate="2009-01-01" firstname="Michael" gender="M" lastname="Pfütsch" license="409144"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="10" heatid="149" lane="1" points="369" resultid="1122" swimtime="00:00:29.13"><SPLITS/></RESULT><RESULT eventid="14" heatid="221" lane="3" points="286" resultid="1676" swimtime="00:01:18.28"><SPLITS><SPLIT distance="50" swimtime="00:00:37.61"/></SPLITS></RESULT><RESULT eventid="28" heatid="284" lane="3" points="305" resultid="2111" swimtime="00:00:35.19"><SPLITS/></RESULT><RESULT eventid="30" heatid="320" lane="4" points="328" resultid="2385" swimtime="00:02:27.78"><SPLITS><SPLIT distance="50" swimtime="00:00:32.11"/><SPLIT distance="100" swimtime="00:01:11.72"/><SPLIT distance="150" swimtime="00:01:51.70"/></SPLITS></RESULT><RESULT eventid="36" heatid="394" lane="5" points="332" resultid="2938" swimtime="00:00:32.13"><SPLITS/></RESULT><RESULT eventid="40" heatid="469" lane="2" points="412" resultid="3507" swimtime="00:01:02.97"><SPLITS><SPLIT distance="50" swimtime="00:00:29.84"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="552" birthdate="2010-01-01" firstname="Noah Nicholas" gender="M" lastname="Murgu" license="436708"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="10" heatid="149" lane="2" points="392" resultid="1123" swimtime="00:00:28.55"><SPLITS/></RESULT><RESULT eventid="14" heatid="223" lane="2" points="352" resultid="1691" swimtime="00:01:13.04"><SPLITS/></RESULT><RESULT eventid="28" heatid="285" lane="6" points="389" resultid="2121" swimtime="00:00:32.46"><SPLITS/></RESULT><RESULT eventid="30" heatid="321" lane="4" points="367" resultid="2391" swimtime="00:02:22.41"><SPLITS><SPLIT distance="50" swimtime="00:00:30.33"/><SPLIT distance="100" swimtime="00:01:06.16"/><SPLIT distance="150" swimtime="00:01:45.28"/></SPLITS></RESULT><RESULT eventid="36" heatid="393" lane="4" points="306" resultid="2929" swimtime="00:00:33.02"><SPLITS/></RESULT><RESULT eventid="40" heatid="469" lane="3" points="410" resultid="3508" swimtime="00:01:03.07"><SPLITS><SPLIT distance="50" swimtime="00:00:29.65"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="553" birthdate="2009-01-01" firstname="Alois" gender="M" lastname="Purbojo" license="409146"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="10" heatid="149" lane="4" points="395" resultid="1125" swimtime="00:00:28.48"><SPLITS/></RESULT><RESULT eventid="12" heatid="182" lane="5" points="301" resultid="1378" swimtime="00:02:49.99"><SPLITS><SPLIT distance="50" swimtime="00:00:34.85"/><SPLIT distance="100" swimtime="00:01:16.90"/><SPLIT distance="150" swimtime="00:02:11.19"/></SPLITS></RESULT><RESULT eventid="28" heatid="284" lane="8" points="280" resultid="2115" swimtime="00:00:36.21"><SPLITS/></RESULT><RESULT eventid="30" heatid="319" lane="3" points="330" resultid="2376" swimtime="00:02:27.58"><SPLITS><SPLIT distance="50" swimtime="00:00:32.35"/><SPLIT distance="100" swimtime="00:01:08.70"/><SPLIT distance="150" swimtime="00:01:47.85"/></SPLITS></RESULT><RESULT eventid="36" heatid="392" lane="2" points="290" resultid="2919" swimtime="00:00:33.62"><SPLITS/></RESULT><RESULT eventid="40" heatid="467" lane="6" points="387" resultid="3495" swimtime="00:01:04.29"><SPLITS><SPLIT distance="50" swimtime="00:00:29.99"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="554" birthdate="2000-01-01" firstname="Maximilian" gender="M" lastname="Ley" license="255969"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="10" heatid="151" lane="8" points="342" resultid="1145" swimtime="00:00:29.89"><SPLITS/></RESULT><RESULT eventid="12" heatid="185" lane="3" points="302" resultid="1398" swimtime="00:02:49.76"><SPLITS><SPLIT distance="50" swimtime="00:00:40.00"/><SPLIT distance="100" swimtime="00:01:21.99"/><SPLIT distance="150" swimtime="00:02:12.92"/></SPLITS></RESULT><RESULT eventid="14" heatid="221" lane="4" points="282" resultid="1677" swimtime="00:01:18.67"><SPLITS><SPLIT distance="50" swimtime="00:00:39.10"/></SPLITS></RESULT><RESULT eventid="32" heatid="354" lane="1" points="301" resultid="2635" swimtime="00:01:24.79"><SPLITS><SPLIT distance="50" swimtime="00:00:40.39"/></SPLITS></RESULT><RESULT eventid="40" heatid="468" lane="6" points="354" resultid="3503" swimtime="00:01:06.18"><SPLITS><SPLIT distance="50" swimtime="00:00:31.40"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="555" birthdate="2007-01-01" firstname="Anton" gender="M" lastname="Grießinger" license="362946"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="10" heatid="153" lane="6" points="466" resultid="1159" swimtime="00:00:26.96"><SPLITS/></RESULT><RESULT eventid="12" heatid="187" lane="4" points="413" resultid="1415" swimtime="00:02:33.06"><SPLITS><SPLIT distance="50" swimtime="00:00:31.47"/><SPLIT distance="100" swimtime="00:01:11.67"/><SPLIT distance="150" swimtime="00:01:59.74"/></SPLITS></RESULT><RESULT eventid="28" heatid="285" lane="5" points="371" resultid="2120" swimtime="00:00:32.98"><SPLITS/></RESULT><RESULT eventid="36" heatid="398" lane="1" points="378" resultid="2966" swimtime="00:00:30.78"><SPLITS/></RESULT><RESULT eventid="40" heatid="474" lane="1" points="454" resultid="3545" swimtime="00:01:00.96"><SPLITS><SPLIT distance="50" swimtime="00:00:28.24"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="571" birthdate="2013-01-01" firstname="Lola" gender="F" lastname="Wening" license="488568"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="27" heatid="254" lane="2" points="99" resultid="1877" swimtime="00:00:58.23"><SPLITS/></RESULT><RESULT eventid="31" heatid="328" lane="3" points="188" resultid="2437" swimtime="00:01:51.83"><SPLITS><SPLIT distance="50" swimtime="00:00:55.86"/></SPLITS></RESULT><RESULT eventid="39" heatid="425" lane="2" points="117" resultid="3164" swimtime="00:01:45.58"><SPLITS><SPLIT distance="50" swimtime="00:00:48.56"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="574" birthdate="2014-01-01" firstname="Victoria" gender="F" lastname="Büttner" license="463010"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="27" heatid="255" lane="2" points="125" resultid="1885" swimtime="00:00:53.82"><SPLITS/></RESULT><RESULT eventid="29" heatid="289" lane="6" points="145" resultid="2148" swimtime="00:03:34.76"><SPLITS><SPLIT distance="50" swimtime="00:00:47.67"/><SPLIT distance="100" swimtime="00:01:43.90"/><SPLIT distance="150" swimtime="00:02:43.78"/></SPLITS></RESULT><RESULT eventid="31" heatid="329" lane="6" points="164" resultid="2448" swimtime="00:01:57.15"><SPLITS><SPLIT distance="50" swimtime="00:00:55.07"/></SPLITS></RESULT><RESULT eventid="39" heatid="424" lane="2" points="151" resultid="3156" swimtime="00:01:37.07"><SPLITS><SPLIT distance="50" swimtime="00:00:46.36"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="575" birthdate="2013-01-01" firstname="Linda" gender="F" lastname="Brand" license="460133"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="27" heatid="256" lane="5" points="162" resultid="1896" swimtime="00:00:49.40"><SPLITS/></RESULT><RESULT eventid="31" heatid="330" lane="6" points="190" resultid="2456" swimtime="00:01:51.50"><SPLITS/></RESULT><RESULT eventid="39" heatid="424" lane="5" points="174" resultid="3159" swimtime="00:01:32.50"><SPLITS><SPLIT distance="50" swimtime="00:00:45.79"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="580" birthdate="2013-01-01" firstname="Laura" gender="F" lastname="Bender" license="462909"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="27" heatid="260" lane="3" points="222" resultid="1926" swimtime="00:00:44.51"><SPLITS/></RESULT><RESULT comment="12:03 Start vor dem Startsignal" eventid="31" heatid="330" lane="7" resultid="2457" status="DSQ" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="39" heatid="425" lane="1" points="220" resultid="3163" swimtime="00:01:25.64"><SPLITS><SPLIT distance="50" swimtime="00:00:40.35"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="582" birthdate="2009-01-01" firstname="Magda" gender="F" lastname="Offinger" license="423316"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="27" heatid="264" lane="3" points="324" resultid="1958" swimtime="00:00:39.26"><SPLITS/></RESULT><RESULT eventid="35" heatid="374" lane="8" points="270" resultid="2789" swimtime="00:00:37.78"><SPLITS/></RESULT><RESULT eventid="39" heatid="437" lane="7" points="293" resultid="3264" swimtime="00:01:17.77"><SPLITS><SPLIT distance="50" swimtime="00:00:36.62"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="586" birthdate="2009-01-01" firstname="Emilia" gender="F" lastname="Kühne" license="404982"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="27" heatid="265" lane="2" points="312" resultid="1965" swimtime="00:00:39.75"><SPLITS/></RESULT><RESULT eventid="29" heatid="300" lane="1" points="293" resultid="2230" swimtime="00:02:49.97"><SPLITS><SPLIT distance="50" swimtime="00:00:37.54"/><SPLIT distance="100" swimtime="00:01:19.06"/><SPLIT distance="150" swimtime="00:02:06.44"/></SPLITS></RESULT><RESULT eventid="35" heatid="372" lane="2" points="247" resultid="2768" swimtime="00:00:38.93"><SPLITS/></RESULT><RESULT eventid="39" heatid="439" lane="5" points="330" resultid="3278" swimtime="00:01:14.78"><SPLITS><SPLIT distance="50" swimtime="00:00:34.95"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="593" birthdate="2011-01-01" firstname="Arno" gender="M" lastname="Lahner" license="455992"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="28" heatid="278" lane="4" points="132" resultid="2064" swimtime="00:00:46.50"><SPLITS/></RESULT><RESULT eventid="30" heatid="311" lane="2" points="136" resultid="2313" swimtime="00:03:18.18"><SPLITS><SPLIT distance="50" swimtime="00:00:42.47"/><SPLIT distance="100" swimtime="00:01:33.44"/><SPLIT distance="150" swimtime="00:02:29.22"/></SPLITS></RESULT><RESULT eventid="40" heatid="456" lane="3" points="132" resultid="3408" swimtime="00:01:31.84"><SPLITS><SPLIT distance="50" swimtime="00:00:43.64"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="609" birthdate="1982-01-01" firstname="André" gender="M" lastname="Kiessg" license="498529"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="36" heatid="390" lane="2" points="201" resultid="2903" swimtime="00:00:37.97"><SPLITS/></RESULT></RESULTS></ATHLETE></ATHLETES><RELAYS><RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="1. Mannschaft" number="1"><ENTRIES/><RESULTS><RESULT eventid="43" heatid="482" lane="3" points="637" resultid="3597" swimtime="00:08:53.73"><SPLITS><SPLIT distance="50" swimtime="00:00:30.33"/><SPLIT distance="100" swimtime="00:01:04.28"/><SPLIT distance="150" swimtime="00:01:39.50"/><SPLIT distance="200" swimtime="00:02:14.06"/><SPLIT distance="250" swimtime="00:02:44.76"/><SPLIT distance="300" swimtime="00:03:18.58"/><SPLIT distance="350" swimtime="00:03:53.54"/><SPLIT distance="400" swimtime="00:04:27.91"/><SPLIT distance="450" swimtime="00:04:59.21"/><SPLIT distance="500" swimtime="00:05:32.41"/><SPLIT distance="550" swimtime="00:06:06.95"/><SPLIT distance="600" swimtime="00:06:40.66"/><SPLIT distance="650" swimtime="00:07:11.23"/><SPLIT distance="700" swimtime="00:07:45.20"/><SPLIT distance="750" swimtime="00:08:20.25"/></SPLITS><RELAYPOSITIONS><RELAYPOSITION athleteid="374" number="1"/><RELAYPOSITION athleteid="179" number="2"/><RELAYPOSITION athleteid="373" number="3"/><RELAYPOSITION athleteid="175" number="4"/></RELAYPOSITIONS></RESULT></RESULTS></RELAY></RELAYS></CLUB><CLUB code="4384" name="SV Wacker Burghausen" nation="GER" region="02" shortname="Burghn" type="CLUB"><CONTACT city="Haag" country="GER" email="svwacker@cmwoods.com" name="Woods, Margarita" phone="017621119729" street="Pfarrer-Kaiser-Ring 34" zip="83527"/><OFFICIALS/><ATHLETES><ATHLETE athleteid="16" birthdate="2017-01-01" firstname="Laura" gender="F" lastname="Verebi" license="483295"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="3" lane="4" points="115" resultid="16" swimtime="00:01:00.20"><SPLITS/></RESULT><RESULT eventid="9" heatid="104" lane="6" points="116" resultid="782" swimtime="00:00:48.46"><SPLITS/></RESULT><RESULT eventid="13" heatid="190" lane="5" points="106" resultid="1438" swimtime="00:02:01.24"><SPLITS/></RESULT><RESULT eventid="27" heatid="254" lane="6" points="116" resultid="1881" swimtime="00:00:55.23"><SPLITS/></RESULT><RESULT eventid="39" heatid="421" lane="7" points="100" resultid="3137" swimtime="00:01:51.29"><SPLITS><SPLIT distance="50" swimtime="00:00:51.46"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="341" birthdate="2013-01-01" firstname="Carolin" gender="F" lastname="Wittig" license="434734"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="47" lane="5" points="429" resultid="356" swimtime="00:05:13.38"><SPLITS><SPLIT distance="100" swimtime="00:01:15.26"/><SPLIT distance="200" swimtime="00:02:36.38"/><SPLIT distance="300" swimtime="00:03:57.19"/></SPLITS></RESULT><RESULT eventid="7" heatid="90" lane="7" points="430" resultid="679" swimtime="00:03:04.07"><SPLITS><SPLIT distance="50" swimtime="00:00:42.07"/><SPLIT distance="100" swimtime="00:01:30.36"/><SPLIT distance="150" swimtime="00:02:18.36"/></SPLITS></RESULT><RESULT eventid="11" heatid="170" lane="7" points="469" resultid="1289" swimtime="00:02:42.30"><SPLITS><SPLIT distance="50" swimtime="00:00:35.10"/><SPLIT distance="100" swimtime="00:01:17.62"/><SPLIT distance="150" swimtime="00:02:05.56"/></SPLITS></RESULT><RESULT eventid="19" heatid="234" lane="5" resultid="1761" swimtime="00:00:52.59"><SPLITS/></RESULT><RESULT eventid="25" heatid="248" lane="7" resultid="1843" swimtime="00:00:50.31"><SPLITS/></RESULT><RESULT eventid="31" heatid="341" lane="3" points="403" resultid="2541" swimtime="00:01:26.82"><SPLITS><SPLIT distance="50" swimtime="00:00:42.00"/></SPLITS></RESULT><RESULT eventid="37" heatid="410" lane="6" points="435" resultid="3060" swimtime="00:02:42.75"><SPLITS><SPLIT distance="50" swimtime="00:00:38.72"/><SPLIT distance="100" swimtime="00:01:20.80"/><SPLIT distance="150" swimtime="00:02:02.55"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="348" birthdate="2012-01-01" firstname="Alina" gender="F" lastname="Iwan" license="404456"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="48" lane="7" points="375" resultid="365" swimtime="00:05:27.70"><SPLITS><SPLIT distance="100" swimtime="00:01:14.03"/><SPLIT distance="200" swimtime="00:02:38.80"/><SPLIT distance="300" swimtime="00:04:05.13"/></SPLITS></RESULT><RESULT eventid="9" heatid="124" lane="4" points="473" resultid="939" swimtime="00:00:30.36"><SPLITS/></RESULT><RESULT eventid="17" heatid="231" lane="8" points="384" resultid="1747" swimtime="00:11:06.61"><SPLITS><SPLIT distance="100" swimtime="00:01:15.34"/><SPLIT distance="200" swimtime="00:02:38.92"/><SPLIT distance="300" swimtime="00:04:04.02"/><SPLIT distance="400" swimtime="00:05:28.95"/><SPLIT distance="500" swimtime="00:06:53.67"/><SPLIT distance="600" swimtime="00:08:19.37"/><SPLIT distance="700" swimtime="00:09:44.80"/></SPLITS></RESULT><RESULT eventid="27" heatid="268" lane="8" points="340" resultid="1995" swimtime="00:00:38.62"><SPLITS/></RESULT><RESULT eventid="29" heatid="302" lane="6" points="431" resultid="2250" swimtime="00:02:29.55"><SPLITS><SPLIT distance="50" swimtime="00:00:33.79"/><SPLIT distance="100" swimtime="00:01:12.66"/><SPLIT distance="150" swimtime="00:01:52.33"/></SPLITS></RESULT><RESULT eventid="35" heatid="372" lane="8" points="315" resultid="2774" swimtime="00:00:35.88"><SPLITS/></RESULT><RESULT eventid="39" heatid="442" lane="5" points="355" resultid="3301" swimtime="00:01:13.01"><SPLITS><SPLIT distance="50" swimtime="00:00:34.45"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="367" birthdate="2011-01-01" firstname="Valentina" gender="F" lastname="Niedermeier" license="417043"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="51" lane="5" points="471" resultid="386" swimtime="00:05:03.78"><SPLITS><SPLIT distance="100" swimtime="00:01:10.65"/><SPLIT distance="200" swimtime="00:02:28.40"/><SPLIT distance="300" swimtime="00:03:46.72"/></SPLITS></RESULT><RESULT eventid="11" heatid="172" lane="5" points="466" resultid="1303" swimtime="00:02:42.62"><SPLITS><SPLIT distance="50" swimtime="00:00:34.99"/><SPLIT distance="100" swimtime="00:01:18.08"/><SPLIT distance="150" swimtime="00:02:06.68"/></SPLITS></RESULT><RESULT eventid="29" heatid="305" lane="3" points="470" resultid="2270" swimtime="00:02:25.25"><SPLITS><SPLIT distance="50" swimtime="00:00:33.58"/><SPLIT distance="100" swimtime="00:01:09.29"/><SPLIT distance="150" swimtime="00:01:48.01"/></SPLITS></RESULT><RESULT eventid="39" heatid="446" lane="5" points="447" resultid="3332" swimtime="00:01:07.58"><SPLITS><SPLIT distance="50" swimtime="00:00:32.33"/></SPLITS></RESULT><RESULT eventid="41" heatid="477" lane="4" points="454" resultid="3566" swimtime="00:05:46.50"><SPLITS><SPLIT distance="50" swimtime="00:00:37.54"/><SPLIT distance="100" swimtime="00:01:22.48"/><SPLIT distance="150" swimtime="00:02:08.62"/><SPLIT distance="200" swimtime="00:02:52.39"/><SPLIT distance="250" swimtime="00:03:42.23"/><SPLIT distance="300" swimtime="00:04:32.08"/><SPLIT distance="350" swimtime="00:05:09.62"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="389" birthdate="2015-01-01" firstname="Theo" gender="M" lastname="Erler" license="464614"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="55" lane="3" points="202" resultid="412" swimtime="00:06:14.48"><SPLITS><SPLIT distance="100" swimtime="00:01:29.73"/><SPLIT distance="200" swimtime="00:03:07.16"/><SPLIT distance="300" swimtime="00:04:43.09"/></SPLITS></RESULT><RESULT eventid="12" heatid="179" lane="8" points="199" resultid="1357" swimtime="00:03:15.01"><SPLITS><SPLIT distance="50" swimtime="00:00:44.49"/><SPLIT distance="100" swimtime="00:01:34.23"/><SPLIT distance="150" swimtime="00:02:31.26"/></SPLITS></RESULT><RESULT eventid="14" heatid="219" lane="8" points="180" resultid="1666" swimtime="00:01:31.33"><SPLITS><SPLIT distance="50" swimtime="00:00:45.58"/></SPLITS></RESULT><RESULT eventid="30" heatid="314" lane="5" points="207" resultid="2338" swimtime="00:02:52.23"><SPLITS><SPLIT distance="50" swimtime="00:00:39.48"/><SPLIT distance="100" swimtime="00:01:25.24"/><SPLIT distance="150" swimtime="00:02:10.15"/></SPLITS></RESULT><RESULT eventid="32" heatid="350" lane="6" points="158" resultid="2609" swimtime="00:01:45.21"><SPLITS><SPLIT distance="50" swimtime="00:00:49.86"/></SPLITS></RESULT><RESULT eventid="36" heatid="388" lane="7" points="139" resultid="2892" swimtime="00:00:42.96"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="432" birthdate="2011-01-01" firstname="Adam" gender="M" lastname="Verebi" license="424450"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="61" lane="7" points="443" resultid="461" swimtime="00:04:48.50"><SPLITS><SPLIT distance="100" swimtime="00:01:10.39"/><SPLIT distance="200" swimtime="00:02:25.05"/><SPLIT distance="300" swimtime="00:03:38.99"/></SPLITS></RESULT><RESULT eventid="6" heatid="78" lane="7" points="389" resultid="588" swimtime="00:01:07.74"><SPLITS><SPLIT distance="50" swimtime="00:00:30.90"/></SPLITS></RESULT><RESULT eventid="10" heatid="152" lane="8" points="410" resultid="1153" swimtime="00:00:28.13"><SPLITS/></RESULT><RESULT eventid="30" heatid="323" lane="6" points="476" resultid="2408" swimtime="00:02:10.57"><SPLITS><SPLIT distance="50" swimtime="00:00:29.83"/><SPLIT distance="100" swimtime="00:01:03.29"/><SPLIT distance="150" swimtime="00:01:37.34"/></SPLITS></RESULT><RESULT eventid="34" heatid="362" lane="1" points="337" resultid="2689" swimtime="00:02:38.45"><SPLITS><SPLIT distance="50" swimtime="00:00:34.69"/><SPLIT distance="100" swimtime="00:01:14.15"/><SPLIT distance="150" swimtime="00:01:56.10"/></SPLITS></RESULT><RESULT eventid="36" heatid="396" lane="7" points="421" resultid="2956" swimtime="00:00:29.70"><SPLITS/></RESULT><RESULT eventid="40" heatid="472" lane="1" points="478" resultid="3530" swimtime="00:00:59.90"><SPLITS><SPLIT distance="50" swimtime="00:00:29.26"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="433" birthdate="2009-01-01" firstname="Daniel" gender="M" lastname="Verebi" license="397410"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="62" lane="1" points="543" resultid="462" swimtime="00:04:29.69"><SPLITS><SPLIT distance="100" swimtime="00:01:01.81"/><SPLIT distance="200" swimtime="00:02:10.06"/><SPLIT distance="300" swimtime="00:03:20.75"/></SPLITS></RESULT><RESULT eventid="10" heatid="154" lane="3" points="454" resultid="1164" swimtime="00:00:27.20"><SPLITS/></RESULT><RESULT eventid="14" heatid="224" lane="4" points="383" resultid="1700" swimtime="00:01:11.03"><SPLITS><SPLIT distance="50" swimtime="00:00:33.20"/></SPLITS></RESULT><RESULT eventid="18" heatid="233" lane="6" points="560" resultid="1757" swimtime="00:09:08.28"><SPLITS><SPLIT distance="100" swimtime="00:01:03.85"/><SPLIT distance="200" swimtime="00:02:12.27"/><SPLIT distance="300" swimtime="00:03:20.20"/><SPLIT distance="400" swimtime="00:04:29.09"/><SPLIT distance="500" swimtime="00:05:38.68"/><SPLIT distance="600" swimtime="00:06:48.99"/><SPLIT distance="700" swimtime="00:07:59.93"/></SPLITS></RESULT><RESULT eventid="30" heatid="324" lane="3" points="536" resultid="2413" swimtime="00:02:05.52"><SPLITS><SPLIT distance="50" swimtime="00:00:28.39"/><SPLIT distance="100" swimtime="00:00:59.70"/><SPLIT distance="150" swimtime="00:01:32.81"/></SPLITS></RESULT><RESULT eventid="36" heatid="396" lane="4" points="419" resultid="2953" swimtime="00:00:29.75"><SPLITS/></RESULT><RESULT eventid="40" heatid="472" lane="6" points="508" resultid="3535" swimtime="00:00:58.71"><SPLITS><SPLIT distance="50" swimtime="00:00:28.09"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="505" birthdate="2009-01-01" firstname="Lennart" gender="M" lastname="Roth" license="406697"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="6" heatid="80" lane="8" points="498" resultid="604" swimtime="00:01:02.36"><SPLITS><SPLIT distance="50" swimtime="00:00:29.11"/></SPLITS></RESULT><RESULT eventid="10" heatid="155" lane="1" points="511" resultid="1169" swimtime="00:00:26.14"><SPLITS/></RESULT><RESULT eventid="34" heatid="362" lane="3" points="374" resultid="2691" swimtime="00:02:33.06"><SPLITS><SPLIT distance="50" swimtime="00:00:31.89"/><SPLIT distance="100" swimtime="00:01:09.71"/><SPLIT distance="150" swimtime="00:01:51.12"/></SPLITS></RESULT><RESULT eventid="36" heatid="399" lane="3" points="506" resultid="2976" swimtime="00:00:27.94"><SPLITS/></RESULT><RESULT eventid="40" heatid="474" lane="5" points="536" resultid="3549" swimtime="00:00:57.68"><SPLITS><SPLIT distance="50" swimtime="00:00:27.59"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="507" birthdate="2012-01-01" firstname="Kassandra" gender="F" lastname="Strohmaier" license="427336"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="7" heatid="91" lane="1" points="481" resultid="681" swimtime="00:02:57.31"><SPLITS><SPLIT distance="50" swimtime="00:00:41.31"/><SPLIT distance="100" swimtime="00:01:27.69"/><SPLIT distance="150" swimtime="00:02:13.60"/></SPLITS></RESULT><RESULT eventid="11" heatid="172" lane="1" points="456" resultid="1299" swimtime="00:02:43.84"><SPLITS><SPLIT distance="50" swimtime="00:00:38.58"/><SPLIT distance="100" swimtime="00:01:20.24"/><SPLIT distance="150" swimtime="00:02:06.57"/></SPLITS></RESULT><RESULT eventid="13" heatid="205" lane="7" points="387" resultid="1558" swimtime="00:01:18.83"><SPLITS><SPLIT distance="50" swimtime="00:00:38.16"/></SPLITS></RESULT><RESULT eventid="31" heatid="343" lane="7" points="462" resultid="2561" swimtime="00:01:22.95"><SPLITS><SPLIT distance="50" swimtime="00:00:39.10"/></SPLITS></RESULT><RESULT eventid="35" heatid="377" lane="8" points="311" resultid="2811" swimtime="00:00:36.02"><SPLITS/></RESULT><RESULT eventid="37" heatid="411" lane="7" points="419" resultid="3069" swimtime="00:02:44.78"><SPLITS><SPLIT distance="100" swimtime="00:01:21.42"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="512" birthdate="2008-01-01" firstname="Tristan" gender="M" lastname="Niedermeier" license="362447"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="8" heatid="101" lane="6" points="474" resultid="761" swimtime="00:02:41.52"><SPLITS><SPLIT distance="50" swimtime="00:00:35.22"/><SPLIT distance="100" swimtime="00:01:17.21"/><SPLIT distance="150" swimtime="00:01:59.15"/></SPLITS></RESULT><RESULT eventid="10" heatid="157" lane="1" points="497" resultid="1184" swimtime="00:00:26.39"><SPLITS/></RESULT><RESULT eventid="32" heatid="356" lane="3" points="461" resultid="2652" swimtime="00:01:13.63"><SPLITS><SPLIT distance="50" swimtime="00:00:34.30"/></SPLITS></RESULT><RESULT eventid="36" heatid="400" lane="7" points="506" resultid="2987" swimtime="00:00:27.93"><SPLITS/></RESULT><RESULT eventid="40" heatid="475" lane="2" points="565" resultid="3553" swimtime="00:00:56.66"><SPLITS><SPLIT distance="50" swimtime="00:00:27.05"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="565" birthdate="2010-01-01" firstname="Hektor" gender="M" lastname="Strohmaier" license="427335"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="12" heatid="188" lane="2" points="462" resultid="1421" swimtime="00:02:27.42"><SPLITS><SPLIT distance="50" swimtime="00:00:31.20"/><SPLIT distance="100" swimtime="00:01:09.14"/><SPLIT distance="150" swimtime="00:01:53.11"/></SPLITS></RESULT><RESULT eventid="14" heatid="224" lane="3" points="445" resultid="1699" swimtime="00:01:07.58"><SPLITS><SPLIT distance="50" swimtime="00:00:32.75"/></SPLITS></RESULT><RESULT eventid="28" heatid="286" lane="5" points="447" resultid="2128" swimtime="00:00:31.00"><SPLITS/></RESULT><RESULT eventid="36" heatid="396" lane="1" points="401" resultid="2950" swimtime="00:00:30.19"><SPLITS/></RESULT><RESULT eventid="38" heatid="419" lane="7" points="446" resultid="3125" swimtime="00:02:26.38"><SPLITS><SPLIT distance="50" swimtime="00:00:33.63"/><SPLIT distance="100" swimtime="00:01:11.33"/><SPLIT distance="150" swimtime="00:01:48.98"/></SPLITS></RESULT><RESULT eventid="40" heatid="471" lane="1" points="458" resultid="3522" swimtime="00:01:00.78"><SPLITS><SPLIT distance="50" swimtime="00:00:29.11"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="608" birthdate="2011-01-01" firstname="Anna" gender="F" lastname="Woods" license="444309"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="35" heatid="379" lane="7" points="362" resultid="2826" swimtime="00:00:34.25"><SPLITS/></RESULT><RESULT eventid="37" heatid="410" lane="4" points="413" resultid="3058" swimtime="00:02:45.59"><SPLITS><SPLIT distance="50" swimtime="00:00:40.18"/><SPLIT distance="100" swimtime="00:01:21.78"/><SPLIT distance="150" swimtime="00:02:03.96"/></SPLITS></RESULT><RESULT eventid="39" heatid="448" lane="2" points="495" resultid="3344" swimtime="00:01:05.34"><SPLITS><SPLIT distance="50" swimtime="00:00:31.34"/></SPLITS></RESULT><RESULT eventid="41" heatid="477" lane="3" points="455" resultid="3565" swimtime="00:05:46.25"><SPLITS><SPLIT distance="50" swimtime="00:00:36.93"/><SPLIT distance="100" swimtime="00:01:19.54"/><SPLIT distance="150" swimtime="00:02:05.20"/><SPLIT distance="200" swimtime="00:02:47.35"/><SPLIT distance="250" swimtime="00:03:40.17"/><SPLIT distance="300" swimtime="00:04:31.47"/><SPLIT distance="350" swimtime="00:05:10.72"/></SPLITS></RESULT></RESULTS></ATHLETE></ATHLETES><RELAYS/></CLUB><CLUB code="4581" name="VSC Donauwörth" nation="GER" region="02" shortname="Donauwör" type="CLUB"><CONTACT city="Donauwörth" country="GER" email="stefanieknab@web.de" name="Lang, Stefanie" phone="0906/20634013" street="Am Zollfeld 4" zip="86609"/><OFFICIALS/><ATHLETES><ATHLETE athleteid="20" birthdate="2017-01-01" firstname="Mathilda" gender="F" lastname="Hauser" license="481461"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="3" lane="8" points="55" resultid="20" swimtime="00:01:16.64"><SPLITS/></RESULT><RESULT eventid="9" heatid="104" lane="1" points="71" resultid="777" swimtime="00:00:56.90"><SPLITS/></RESULT><RESULT eventid="13" heatid="190" lane="3" points="55" resultid="1436" swimtime="00:02:30.18"><SPLITS><SPLIT distance="50" swimtime="00:01:12.51"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="342" birthdate="2011-01-01" firstname="Dora" gender="F" lastname="Pajtas" license="421964"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="47" lane="6" points="343" resultid="357" swimtime="00:05:37.55"><SPLITS><SPLIT distance="100" swimtime="00:01:25.28"/><SPLIT distance="200" swimtime="00:02:41.75"/><SPLIT distance="300" swimtime="00:04:10.37"/></SPLITS></RESULT><RESULT eventid="9" heatid="124" lane="7" points="431" resultid="942" swimtime="00:00:31.32"><SPLITS/></RESULT><RESULT eventid="13" heatid="207" lane="6" points="407" resultid="1572" swimtime="00:01:17.46"><SPLITS><SPLIT distance="50" swimtime="00:00:37.22"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="354" birthdate="2013-01-01" firstname="Elena" gender="F" lastname="Hauser" license="458548"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="49" lane="5" points="436" resultid="371" swimtime="00:05:11.74"><SPLITS><SPLIT distance="100" swimtime="00:01:13.53"/><SPLIT distance="200" swimtime="00:02:33.57"/><SPLIT distance="300" swimtime="00:03:54.24"/></SPLITS></RESULT><RESULT eventid="5" heatid="68" lane="8" points="328" resultid="511" swimtime="00:01:20.37"><SPLITS><SPLIT distance="50" swimtime="00:00:36.96"/></SPLITS></RESULT><RESULT eventid="11" heatid="171" lane="5" points="445" resultid="1295" swimtime="00:02:45.17"><SPLITS><SPLIT distance="50" swimtime="00:00:35.96"/><SPLIT distance="100" swimtime="00:01:18.98"/><SPLIT distance="150" swimtime="00:02:07.44"/></SPLITS></RESULT><RESULT eventid="13" heatid="207" lane="7" points="363" resultid="1573" swimtime="00:01:20.47"><SPLITS><SPLIT distance="50" swimtime="00:00:38.01"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="410" birthdate="2012-01-01" firstname="Moritz" gender="M" lastname="Lang" license="406618"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="58" lane="6" points="336" resultid="439" swimtime="00:05:16.53"><SPLITS><SPLIT distance="100" swimtime="00:01:13.59"/><SPLIT distance="200" swimtime="00:02:35.09"/><SPLIT distance="300" swimtime="00:03:57.97"/></SPLITS></RESULT><RESULT eventid="6" heatid="74" lane="6" points="198" resultid="556" swimtime="00:01:24.83"><SPLITS><SPLIT distance="50" swimtime="00:00:38.16"/></SPLITS></RESULT><RESULT eventid="12" heatid="184" lane="7" points="293" resultid="1394" swimtime="00:02:51.48"><SPLITS><SPLIT distance="50" swimtime="00:00:38.38"/><SPLIT distance="100" swimtime="00:01:21.33"/><SPLIT distance="150" swimtime="00:02:13.62"/></SPLITS></RESULT><RESULT eventid="14" heatid="221" lane="5" points="268" resultid="1678" swimtime="00:01:19.98"><SPLITS><SPLIT distance="50" swimtime="00:00:39.51"/></SPLITS></RESULT></RESULTS></ATHLETE></ATHLETES><RELAYS/></CLUB><CLUB code="4296" name="SC Wfr. München" nation="GER" region="02" shortname="WfrMünch" type="CLUB"><CONTACT city="München" country="GER" email="meldewesen@scw-muenchen.de" name="Killiches, Matthias" phone="+49 172 8563528" street="Lazarettstraße 5" zip="80636"/><OFFICIALS/><ATHLETES><ATHLETE athleteid="21" birthdate="2016-01-01" firstname="Selma" gender="F" lastname="Burkhart" license="473761"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="4" lane="1" points="101" resultid="21" swimtime="00:01:02.80"><SPLITS/></RESULT><RESULT eventid="9" heatid="104" lane="4" points="159" resultid="780" swimtime="00:00:43.62"><SPLITS/></RESULT><RESULT eventid="13" heatid="193" lane="3" points="126" resultid="1458" swimtime="00:01:54.51"><SPLITS><SPLIT distance="50" swimtime="00:00:57.65"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="42" birthdate="2017-01-01" firstname="Giulia" gender="F" lastname="Spang" license="495524"><HANDICAP/><ENTRIES/><RESULTS><RESULT comment="09:16 Start vor dem Startsignal" eventid="1" heatid="6" lane="6" resultid="42" status="DSQ" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="9" heatid="108" lane="1" points="119" resultid="809" swimtime="00:00:48.01"><SPLITS/></RESULT><RESULT eventid="27" heatid="257" lane="4" points="152" resultid="1903" swimtime="00:00:50.48"><SPLITS/></RESULT><RESULT eventid="39" heatid="422" lane="2" points="103" resultid="3140" swimtime="00:01:49.97"><SPLITS><SPLIT distance="50" swimtime="00:00:50.04"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="60" birthdate="2016-01-01" firstname="Nura" gender="F" lastname="Al-Sultan" license="464789"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="8" lane="8" points="197" resultid="60" swimtime="00:00:50.32"><SPLITS/></RESULT><RESULT eventid="9" heatid="110" lane="1" points="254" resultid="825" swimtime="00:00:37.35"><SPLITS/></RESULT><RESULT eventid="13" heatid="193" lane="4" points="199" resultid="1459" swimtime="00:01:38.24"><SPLITS><SPLIT distance="50" swimtime="00:00:48.45"/></SPLITS></RESULT><RESULT eventid="29" heatid="292" lane="1" points="233" resultid="2166" swimtime="00:03:03.48"><SPLITS><SPLIT distance="50" swimtime="00:00:43.22"/><SPLIT distance="100" swimtime="00:01:31.97"/><SPLIT distance="150" swimtime="00:02:20.16"/></SPLITS></RESULT><RESULT eventid="31" heatid="331" lane="3" points="193" resultid="2461" swimtime="00:01:50.82"><SPLITS/></RESULT><RESULT eventid="39" heatid="429" lane="7" points="213" resultid="3200" swimtime="00:01:26.49"><SPLITS><SPLIT distance="50" swimtime="00:00:40.89"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="65" birthdate="2017-01-01" firstname="Lena" gender="F" lastname="Rauschmayr" license="493646"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="9" lane="5" points="158" resultid="65" swimtime="00:00:54.17"><SPLITS/></RESULT><RESULT eventid="9" heatid="106" lane="2" points="136" resultid="794" swimtime="00:00:45.94"><SPLITS/></RESULT><RESULT eventid="27" heatid="259" lane="7" points="173" resultid="1922" swimtime="00:00:48.36"><SPLITS/></RESULT><RESULT eventid="39" heatid="424" lane="6" points="123" resultid="3160" swimtime="00:01:43.78"><SPLITS><SPLIT distance="50" swimtime="00:00:47.91"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="77" birthdate="2015-01-01" firstname="Sofia" gender="F" lastname="Spang" license="470052"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="11" lane="1" points="198" resultid="77" swimtime="00:00:50.20"><SPLITS/></RESULT><RESULT eventid="5" heatid="63" lane="3" points="140" resultid="469" swimtime="00:01:46.78"><SPLITS><SPLIT distance="50" swimtime="00:00:47.36"/></SPLITS></RESULT><RESULT eventid="13" heatid="195" lane="2" points="213" resultid="1473" swimtime="00:01:36.17"><SPLITS><SPLIT distance="50" swimtime="00:00:47.73"/></SPLITS></RESULT><RESULT eventid="31" heatid="333" lane="8" points="212" resultid="2482" swimtime="00:01:47.45"><SPLITS><SPLIT distance="50" swimtime="00:00:50.70"/></SPLITS></RESULT><RESULT eventid="39" heatid="429" lane="1" points="217" resultid="3194" swimtime="00:01:26.04"><SPLITS><SPLIT distance="50" swimtime="00:00:41.40"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="111" birthdate="2012-01-01" firstname="Eva" gender="F" lastname="Schreiner" license="420331"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="15" lane="3" points="254" resultid="111" swimtime="00:00:46.25"><SPLITS/></RESULT><RESULT eventid="3" heatid="47" lane="3" points="380" resultid="354" swimtime="00:05:26.36"><SPLITS><SPLIT distance="100" swimtime="00:01:16.72"/><SPLIT distance="200" swimtime="00:02:40.28"/><SPLIT distance="300" swimtime="00:04:04.36"/></SPLITS></RESULT><RESULT eventid="9" heatid="119" lane="3" points="342" resultid="898" swimtime="00:00:33.82"><SPLITS/></RESULT><RESULT eventid="13" heatid="202" lane="4" points="321" resultid="1531" swimtime="00:01:23.89"><SPLITS><SPLIT distance="50" swimtime="00:00:40.42"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="121" birthdate="2010-01-01" firstname="Marie-Christin" gender="F" lastname="Karras" license="440553"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="16" lane="5" points="287" resultid="121" swimtime="00:00:44.40"><SPLITS/></RESULT><RESULT eventid="5" heatid="66" lane="3" points="343" resultid="491" swimtime="00:01:19.19"><SPLITS><SPLIT distance="50" swimtime="00:00:35.31"/></SPLITS></RESULT><RESULT eventid="9" heatid="124" lane="1" points="429" resultid="936" swimtime="00:00:31.36"><SPLITS/></RESULT><RESULT eventid="27" heatid="265" lane="5" points="357" resultid="1968" swimtime="00:00:38.01"><SPLITS/></RESULT><RESULT eventid="29" heatid="301" lane="8" points="399" resultid="2244" swimtime="00:02:33.40"><SPLITS><SPLIT distance="50" swimtime="00:00:34.45"/><SPLIT distance="100" swimtime="00:01:13.43"/><SPLIT distance="150" swimtime="00:01:55.37"/></SPLITS></RESULT><RESULT eventid="35" heatid="375" lane="3" points="326" resultid="2792" swimtime="00:00:35.47"><SPLITS/></RESULT><RESULT eventid="39" heatid="441" lane="3" points="422" resultid="3291" swimtime="00:01:08.91"><SPLITS><SPLIT distance="50" swimtime="00:00:33.41"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="127" birthdate="2013-01-01" firstname="Elli" gender="F" lastname="Glashauser" license="453832"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="17" lane="3" points="286" resultid="127" swimtime="00:00:44.45"><SPLITS/></RESULT><RESULT eventid="7" heatid="88" lane="5" points="351" resultid="661" swimtime="00:03:16.82"><SPLITS><SPLIT distance="50" swimtime="00:00:46.02"/><SPLIT distance="100" swimtime="00:01:37.59"/><SPLIT distance="150" swimtime="00:02:28.53"/></SPLITS></RESULT><RESULT eventid="11" heatid="167" lane="5" points="374" resultid="1263" swimtime="00:02:54.92"><SPLITS><SPLIT distance="50" swimtime="00:00:41.05"/><SPLIT distance="100" swimtime="00:01:27.37"/><SPLIT distance="150" swimtime="00:02:16.82"/></SPLITS></RESULT><RESULT eventid="25" heatid="248" lane="5" resultid="1841" swimtime="00:00:55.49"><SPLITS/></RESULT><RESULT eventid="29" heatid="299" lane="2" points="335" resultid="2223" swimtime="00:02:42.67"><SPLITS><SPLIT distance="50" swimtime="00:00:38.48"/><SPLIT distance="100" swimtime="00:01:20.19"/><SPLIT distance="150" swimtime="00:02:03.85"/></SPLITS></RESULT><RESULT eventid="31" heatid="338" lane="3" points="327" resultid="2517" swimtime="00:01:33.07"><SPLITS><SPLIT distance="50" swimtime="00:00:45.72"/></SPLITS></RESULT><RESULT eventid="39" heatid="437" lane="1" points="347" resultid="3258" swimtime="00:01:13.54"><SPLITS><SPLIT distance="50" swimtime="00:00:36.22"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="140" birthdate="2002-01-01" firstname="Hanna" gender="F" lastname="Pretzlik" license="404246"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="18" lane="8" points="306" resultid="140" swimtime="00:00:43.44"><SPLITS/></RESULT><RESULT eventid="7" heatid="88" lane="6" points="334" resultid="662" swimtime="00:03:20.11"><SPLITS><SPLIT distance="50" swimtime="00:00:46.39"/><SPLIT distance="100" swimtime="00:01:37.30"/><SPLIT distance="150" swimtime="00:02:29.70"/></SPLITS></RESULT><RESULT eventid="9" heatid="117" lane="4" points="360" resultid="883" swimtime="00:00:33.26"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="151" birthdate="2012-01-01" firstname="Greta" gender="F" lastname="Glashauser" license="436953"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="20" lane="3" points="410" resultid="151" swimtime="00:00:39.42"><SPLITS/></RESULT><RESULT eventid="7" heatid="90" lane="6" points="437" resultid="678" swimtime="00:03:03.05"><SPLITS><SPLIT distance="50" swimtime="00:00:40.90"/><SPLIT distance="100" swimtime="00:01:28.36"/><SPLIT distance="150" swimtime="00:02:16.22"/></SPLITS></RESULT><RESULT eventid="15" heatid="226" lane="3" points="376" resultid="1714" swimtime="00:21:14.97"><SPLITS><SPLIT distance="100" swimtime="00:01:17.15"/><SPLIT distance="200" swimtime="00:02:41.46"/><SPLIT distance="300" swimtime="00:04:07.28"/><SPLIT distance="400" swimtime="00:05:31.77"/><SPLIT distance="500" swimtime="00:06:56.84"/><SPLIT distance="600" swimtime="00:08:22.55"/><SPLIT distance="700" swimtime="00:09:47.87"/><SPLIT distance="800" swimtime="00:11:13.42"/><SPLIT distance="900" swimtime="00:12:38.86"/><SPLIT distance="1000" swimtime="00:14:04.51"/><SPLIT distance="1100" swimtime="00:15:31.22"/><SPLIT distance="1200" swimtime="00:16:58.07"/><SPLIT distance="1300" swimtime="00:18:24.63"/><SPLIT distance="1400" swimtime="00:19:51.12"/></SPLITS></RESULT><RESULT eventid="31" heatid="341" lane="1" points="430" resultid="2539" swimtime="00:01:24.92"><SPLITS><SPLIT distance="50" swimtime="00:00:40.13"/></SPLITS></RESULT><RESULT eventid="33" heatid="358" lane="5" points="269" resultid="2664" swimtime="00:03:08.66"><SPLITS><SPLIT distance="50" swimtime="00:00:38.89"/><SPLIT distance="100" swimtime="00:01:27.86"/><SPLIT distance="150" swimtime="00:02:19.17"/></SPLITS></RESULT><RESULT eventid="35" heatid="375" lane="7" points="299" resultid="2796" swimtime="00:00:36.51"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="154" birthdate="2012-01-01" firstname="Laetitia" gender="F" lastname="Adelhardt" license="419158"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="20" lane="6" points="408" resultid="154" swimtime="00:00:39.50"><SPLITS/></RESULT><RESULT eventid="5" heatid="70" lane="4" points="523" resultid="523" swimtime="00:01:08.82"><SPLITS><SPLIT distance="50" swimtime="00:00:33.01"/></SPLITS></RESULT><RESULT eventid="11" heatid="173" lane="5" points="524" resultid="1311" swimtime="00:02:36.36"><SPLITS><SPLIT distance="50" swimtime="00:00:33.02"/><SPLIT distance="100" swimtime="00:01:12.41"/><SPLIT distance="150" swimtime="00:02:00.11"/></SPLITS></RESULT><RESULT eventid="13" heatid="209" lane="7" points="561" resultid="1588" swimtime="00:01:09.64"><SPLITS><SPLIT distance="50" swimtime="00:00:34.41"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="168" birthdate="2009-01-01" firstname="Elena" gender="F" lastname="Schreiber" license="414371"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="22" lane="6" points="388" resultid="168" swimtime="00:00:40.17"><SPLITS/></RESULT><RESULT eventid="9" heatid="126" lane="2" points="446" resultid="953" swimtime="00:00:30.96"><SPLITS/></RESULT><RESULT eventid="17" heatid="231" lane="6" points="317" resultid="1745" swimtime="00:11:50.71"><SPLITS><SPLIT distance="100" swimtime="00:01:13.61"/><SPLIT distance="200" swimtime="00:02:39.47"/><SPLIT distance="300" swimtime="00:04:09.78"/><SPLIT distance="400" swimtime="00:05:42.76"/><SPLIT distance="500" swimtime="00:07:16.62"/><SPLIT distance="600" swimtime="00:08:49.81"/><SPLIT distance="700" swimtime="00:10:22.36"/></SPLITS></RESULT><RESULT eventid="27" heatid="269" lane="2" points="417" resultid="1997" swimtime="00:00:36.11"><SPLITS/></RESULT><RESULT eventid="35" heatid="376" lane="7" points="346" resultid="2804" swimtime="00:00:34.78"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="185" birthdate="2011-01-01" firstname="Leonie" gender="F" lastname="Platzer" license="416840"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="24" lane="7" points="533" resultid="185" swimtime="00:00:36.13"><SPLITS/></RESULT><RESULT eventid="9" heatid="129" lane="4" points="498" resultid="978" swimtime="00:00:29.86"><SPLITS/></RESULT><RESULT eventid="29" heatid="305" lane="8" points="505" resultid="2274" swimtime="00:02:21.86"><SPLITS><SPLIT distance="50" swimtime="00:00:32.87"/><SPLIT distance="100" swimtime="00:01:08.17"/><SPLIT distance="150" swimtime="00:01:45.82"/></SPLITS></RESULT><RESULT eventid="31" heatid="342" lane="4" points="439" resultid="2550" swimtime="00:01:24.35"><SPLITS><SPLIT distance="50" swimtime="00:00:39.96"/></SPLITS></RESULT><RESULT eventid="35" heatid="382" lane="2" points="501" resultid="2845" swimtime="00:00:30.74"><SPLITS/></RESULT><RESULT eventid="39" heatid="447" lane="6" points="437" resultid="3340" swimtime="00:01:08.12"><SPLITS><SPLIT distance="50" swimtime="00:00:32.23"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="194" birthdate="2013-01-01" firstname="Lorenzo" gender="M" lastname="Simeone" license="486366"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="26" lane="5" points="120" resultid="194" swimtime="00:00:52.54"><SPLITS/></RESULT><RESULT eventid="10" heatid="134" lane="3" points="127" resultid="1008" swimtime="00:00:41.59"><SPLITS/></RESULT><RESULT eventid="14" heatid="210" lane="2" points="106" resultid="1591" swimtime="00:01:48.96"><SPLITS><SPLIT distance="50" swimtime="00:00:51.62"/></SPLITS></RESULT><RESULT eventid="30" heatid="309" lane="1" points="106" resultid="2296" swimtime="00:03:35.35"><SPLITS><SPLIT distance="50" swimtime="00:00:47.29"/><SPLIT distance="100" swimtime="00:01:41.79"/><SPLIT distance="150" swimtime="00:02:42.54"/></SPLITS></RESULT><RESULT eventid="32" heatid="346" lane="1" points="107" resultid="2575" swimtime="00:01:59.72"><SPLITS><SPLIT distance="50" swimtime="00:00:57.26"/></SPLITS></RESULT><RESULT eventid="36" heatid="384" lane="5" points="68" resultid="2859" swimtime="00:00:54.33"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="204" birthdate="2017-01-01" firstname="Patrik" gender="M" lastname="Csontos" license="500734"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="27" lane="8" points="82" resultid="204" swimtime="00:00:59.68"><SPLITS/></RESULT><RESULT eventid="10" heatid="134" lane="1" points="78" resultid="1006" swimtime="00:00:48.80"><SPLITS/></RESULT><RESULT eventid="28" heatid="274" lane="7" points="86" resultid="2037" swimtime="00:00:53.66"><SPLITS/></RESULT><RESULT eventid="40" heatid="453" lane="8" points="62" resultid="3389" swimtime="00:01:57.81"><SPLITS><SPLIT distance="50" swimtime="00:00:59.27"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="213" birthdate="2014-01-01" firstname="Elias" gender="M" lastname="Schober" license="495935"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="29" lane="1" points="95" resultid="213" swimtime="00:00:56.78"><SPLITS/></RESULT><RESULT eventid="10" heatid="137" lane="2" points="120" resultid="1030" swimtime="00:00:42.37"><SPLITS/></RESULT><RESULT eventid="14" heatid="213" lane="8" points="119" resultid="1620" swimtime="00:01:44.85"><SPLITS><SPLIT distance="50" swimtime="00:00:52.26"/></SPLITS></RESULT><RESULT eventid="28" heatid="278" lane="5" points="117" resultid="2065" swimtime="00:00:48.45"><SPLITS/></RESULT><RESULT eventid="32" heatid="346" lane="4" points="79" resultid="2578" swimtime="00:02:12.36"><SPLITS><SPLIT distance="50" swimtime="00:01:00.24"/></SPLITS></RESULT><RESULT eventid="36" heatid="385" lane="3" points="51" resultid="2865" swimtime="00:00:59.83"><SPLITS/></RESULT><RESULT eventid="40" heatid="456" lane="8" points="111" resultid="3412" swimtime="00:01:37.46"><SPLITS><SPLIT distance="50" swimtime="00:00:45.02"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="216" birthdate="2014-01-01" firstname="Johannes" gender="M" lastname="Nibler" license="451233"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="29" lane="4" points="146" resultid="216" swimtime="00:00:49.21"><SPLITS/></RESULT><RESULT eventid="10" heatid="142" lane="8" points="177" resultid="1074" swimtime="00:00:37.20"><SPLITS/></RESULT><RESULT eventid="12" heatid="177" lane="4" points="186" resultid="1338" swimtime="00:03:19.38"><SPLITS><SPLIT distance="50" swimtime="00:00:42.30"/><SPLIT distance="100" swimtime="00:01:32.73"/><SPLIT distance="150" swimtime="00:02:32.81"/></SPLITS></RESULT><RESULT eventid="30" heatid="314" lane="7" points="193" resultid="2340" swimtime="00:02:56.45"><SPLITS><SPLIT distance="50" swimtime="00:00:38.71"/><SPLIT distance="100" swimtime="00:01:24.66"/><SPLIT distance="150" swimtime="00:02:10.77"/></SPLITS></RESULT><RESULT eventid="36" heatid="389" lane="7" points="141" resultid="2900" swimtime="00:00:42.71"><SPLITS/></RESULT><RESULT eventid="40" heatid="460" lane="1" points="183" resultid="3437" swimtime="00:01:22.44"><SPLITS><SPLIT distance="50" swimtime="00:00:39.14"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="226" birthdate="2014-01-01" firstname="Quirin" gender="M" lastname="Thiele" license="481241"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="30" lane="6" points="139" resultid="226" swimtime="00:00:50.08"><SPLITS/></RESULT><RESULT eventid="4" heatid="53" lane="2" points="166" resultid="398" swimtime="00:06:40.12"><SPLITS><SPLIT distance="100" swimtime="00:01:34.15"/><SPLIT distance="200" swimtime="00:03:18.47"/><SPLIT distance="300" swimtime="00:05:03.97"/></SPLITS></RESULT><RESULT eventid="14" heatid="216" lane="4" points="152" resultid="1638" swimtime="00:01:36.66"><SPLITS><SPLIT distance="50" swimtime="00:00:45.62"/></SPLITS></RESULT><RESULT eventid="26" heatid="250" lane="3" resultid="1853" swimtime="00:01:03.66"><SPLITS/></RESULT><RESULT eventid="32" heatid="348" lane="6" points="143" resultid="2595" swimtime="00:01:48.55"><SPLITS><SPLIT distance="50" swimtime="00:00:52.23"/></SPLITS></RESULT><RESULT eventid="40" heatid="458" lane="6" points="175" resultid="3426" swimtime="00:01:23.70"><SPLITS><SPLIT distance="50" swimtime="00:00:39.81"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="229" birthdate="2015-01-01" firstname="Theodor" gender="M" lastname="Engelmann" license="464839"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="31" lane="1" points="151" resultid="229" swimtime="00:00:48.69"><SPLITS/></RESULT><RESULT eventid="8" heatid="95" lane="1" points="182" resultid="712" swimtime="00:03:42.21"><SPLITS><SPLIT distance="50" swimtime="00:00:52.67"/><SPLIT distance="100" swimtime="00:01:49.82"/><SPLIT distance="150" swimtime="00:02:50.94"/></SPLITS></RESULT><RESULT eventid="14" heatid="217" lane="1" points="180" resultid="1643" swimtime="00:01:31.31"><SPLITS><SPLIT distance="50" swimtime="00:00:46.41"/></SPLITS></RESULT><RESULT eventid="30" heatid="312" lane="8" points="173" resultid="2326" swimtime="00:03:02.73"><SPLITS><SPLIT distance="50" swimtime="00:00:42.33"/><SPLIT distance="100" swimtime="00:01:28.76"/><SPLIT distance="150" swimtime="00:02:17.93"/></SPLITS></RESULT><RESULT eventid="36" heatid="384" lane="3" points="102" resultid="2857" swimtime="00:00:47.65"><SPLITS/></RESULT><RESULT eventid="40" heatid="457" lane="6" points="174" resultid="3418" swimtime="00:01:23.89"><SPLITS><SPLIT distance="50" swimtime="00:00:40.58"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="238" birthdate="2012-01-01" firstname="Simeon" gender="M" lastname="Tokaji" license="433820"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="32" lane="2" points="177" resultid="238" swimtime="00:00:46.14"><SPLITS/></RESULT><RESULT eventid="12" heatid="182" lane="3" points="236" resultid="1376" swimtime="00:03:04.45"><SPLITS><SPLIT distance="50" swimtime="00:00:40.84"/><SPLIT distance="100" swimtime="00:01:27.53"/><SPLIT distance="150" swimtime="00:02:23.92"/></SPLITS></RESULT><RESULT eventid="18" heatid="232" lane="3" resultid="1749" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="30" heatid="319" lane="1" points="278" resultid="2374" swimtime="00:02:36.28"><SPLITS><SPLIT distance="50" swimtime="00:00:37.73"/><SPLIT distance="100" swimtime="00:01:16.36"/><SPLIT distance="150" swimtime="00:01:57.01"/></SPLITS></RESULT><RESULT eventid="32" heatid="350" lane="2" points="179" resultid="2606" swimtime="00:01:40.87"><SPLITS><SPLIT distance="50" swimtime="00:00:49.31"/></SPLITS></RESULT><RESULT eventid="36" heatid="390" lane="5" points="200" resultid="2906" swimtime="00:00:38.08"><SPLITS/></RESULT><RESULT eventid="40" heatid="464" lane="6" points="259" resultid="3472" swimtime="00:01:13.44"><SPLITS><SPLIT distance="50" swimtime="00:00:35.45"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="253" birthdate="2013-01-01" firstname="Jonas" gender="M" lastname="Festerling" license="453165"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="34" lane="1" points="177" resultid="253" swimtime="00:00:46.14"><SPLITS/></RESULT><RESULT eventid="8" heatid="97" lane="1" points="195" resultid="726" swimtime="00:03:37.09"><SPLITS><SPLIT distance="50" swimtime="00:00:49.35"/><SPLIT distance="100" swimtime="00:01:45.28"/><SPLIT distance="150" swimtime="00:02:44.08"/></SPLITS></RESULT><RESULT eventid="12" heatid="179" lane="7" points="225" resultid="1356" swimtime="00:03:07.34"><SPLITS><SPLIT distance="50" swimtime="00:00:44.95"/><SPLIT distance="100" swimtime="00:01:36.64"/><SPLIT distance="150" swimtime="00:02:27.82"/></SPLITS></RESULT><RESULT eventid="30" heatid="317" lane="8" points="234" resultid="2365" swimtime="00:02:45.32"><SPLITS><SPLIT distance="50" swimtime="00:00:37.69"/><SPLIT distance="100" swimtime="00:01:18.80"/><SPLIT distance="150" swimtime="00:02:03.82"/></SPLITS></RESULT><RESULT eventid="32" heatid="350" lane="1" points="183" resultid="2605" swimtime="00:01:40.12"><SPLITS><SPLIT distance="50" swimtime="00:00:50.58"/></SPLITS></RESULT><RESULT eventid="36" heatid="386" lane="8" points="123" resultid="2878" swimtime="00:00:44.74"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="254" birthdate="2011-01-01" firstname="Alexander" gender="M" lastname="Weizel" license="419161"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="34" lane="2" points="182" resultid="254" swimtime="00:00:45.73"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="263" birthdate="2011-01-01" firstname="Henry" gender="M" lastname="Müller" license="416820"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="35" lane="5" points="244" resultid="263" swimtime="00:00:41.51"><SPLITS/></RESULT><RESULT eventid="4" heatid="58" lane="4" points="310" resultid="437" swimtime="00:05:24.82"><SPLITS><SPLIT distance="100" swimtime="00:01:15.05"/><SPLIT distance="200" swimtime="00:02:38.08"/><SPLIT distance="300" swimtime="00:04:02.36"/></SPLITS></RESULT><RESULT eventid="10" heatid="145" lane="7" points="244" resultid="1096" swimtime="00:00:33.42"><SPLITS/></RESULT><RESULT eventid="14" heatid="220" lane="8" points="253" resultid="1673" swimtime="00:01:21.50"><SPLITS><SPLIT distance="50" swimtime="00:00:39.67"/></SPLITS></RESULT><RESULT eventid="28" heatid="282" lane="6" points="258" resultid="2098" swimtime="00:00:37.20"><SPLITS/></RESULT><RESULT eventid="30" heatid="319" lane="7" points="295" resultid="2380" swimtime="00:02:33.16"><SPLITS><SPLIT distance="50" swimtime="00:00:34.83"/><SPLIT distance="100" swimtime="00:01:14.37"/><SPLIT distance="150" swimtime="00:01:54.66"/></SPLITS></RESULT><RESULT eventid="32" heatid="351" lane="4" points="230" resultid="2615" swimtime="00:01:32.75"><SPLITS><SPLIT distance="50" swimtime="00:00:43.62"/></SPLITS></RESULT><RESULT eventid="38" heatid="417" lane="4" points="277" resultid="3110" swimtime="00:02:51.62"><SPLITS><SPLIT distance="50" swimtime="00:00:40.01"/><SPLIT distance="100" swimtime="00:01:24.34"/><SPLIT distance="150" swimtime="00:02:08.63"/></SPLITS></RESULT><RESULT eventid="40" heatid="465" lane="8" points="263" resultid="3482" swimtime="00:01:13.06"><SPLITS><SPLIT distance="50" swimtime="00:00:35.18"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="266" birthdate="2011-01-01" firstname="Alan Julian" gender="M" lastname="Said" license="431637"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="35" lane="8" points="213" resultid="266" swimtime="00:00:43.45"><SPLITS/></RESULT><RESULT eventid="8" heatid="97" lane="5" points="234" resultid="730" swimtime="00:03:24.25"><SPLITS><SPLIT distance="50" swimtime="00:00:46.99"/><SPLIT distance="100" swimtime="00:01:40.00"/><SPLIT distance="150" swimtime="00:02:33.18"/></SPLITS></RESULT><RESULT eventid="10" heatid="144" lane="2" points="236" resultid="1083" swimtime="00:00:33.79"><SPLITS/></RESULT><RESULT eventid="18" heatid="232" lane="2" points="252" resultid="1748" swimtime="00:11:55.25"><SPLITS><SPLIT distance="100" swimtime="00:01:23.63"/><SPLIT distance="200" swimtime="00:02:55.42"/><SPLIT distance="300" swimtime="00:04:26.99"/><SPLIT distance="400" swimtime="00:05:58.74"/><SPLIT distance="500" swimtime="00:07:30.03"/><SPLIT distance="600" swimtime="00:09:01.80"/><SPLIT distance="700" swimtime="00:10:32.16"/></SPLITS></RESULT><RESULT eventid="32" heatid="351" lane="2" points="222" resultid="2613" swimtime="00:01:33.80"><SPLITS><SPLIT distance="50" swimtime="00:00:46.20"/></SPLITS></RESULT><RESULT eventid="38" heatid="416" lane="8" points="236" resultid="3106" swimtime="00:03:00.90"><SPLITS><SPLIT distance="50" swimtime="00:00:44.05"/><SPLIT distance="100" swimtime="00:01:29.41"/><SPLIT distance="150" swimtime="00:02:16.92"/></SPLITS></RESULT><RESULT eventid="40" heatid="462" lane="4" points="231" resultid="3455" swimtime="00:01:16.27"><SPLITS><SPLIT distance="50" swimtime="00:00:35.74"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="281" birthdate="2011-01-01" firstname="Toni" gender="M" lastname="Krizanovic" license="443243"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="37" lane="7" points="343" resultid="281" swimtime="00:00:37.04"><SPLITS/></RESULT><RESULT eventid="8" heatid="100" lane="8" points="326" resultid="756" swimtime="00:03:02.86"><SPLITS><SPLIT distance="50" swimtime="00:00:42.39"/><SPLIT distance="100" swimtime="00:01:28.85"/><SPLIT distance="150" swimtime="00:02:17.55"/></SPLITS></RESULT><RESULT eventid="10" heatid="146" lane="5" points="299" resultid="1102" swimtime="00:00:31.27"><SPLITS/></RESULT><RESULT eventid="12" heatid="181" lane="3" points="299" resultid="1368" swimtime="00:02:50.35"><SPLITS><SPLIT distance="50" swimtime="00:00:38.03"/><SPLIT distance="100" swimtime="00:01:26.58"/><SPLIT distance="150" swimtime="00:02:13.17"/></SPLITS></RESULT><RESULT eventid="32" heatid="353" lane="3" points="334" resultid="2629" swimtime="00:01:21.96"><SPLITS><SPLIT distance="50" swimtime="00:00:39.44"/></SPLITS></RESULT><RESULT eventid="40" heatid="465" lane="4" points="295" resultid="3478" swimtime="00:01:10.38"><SPLITS><SPLIT distance="50" swimtime="00:00:34.54"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="285" birthdate="2010-01-01" firstname="Hugo" gender="M" lastname="Liedl" license="410668"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="38" lane="3" points="397" resultid="285" swimtime="00:00:35.28"><SPLITS/></RESULT><RESULT eventid="8" heatid="98" lane="5" points="414" resultid="737" swimtime="00:02:48.86"><SPLITS><SPLIT distance="50" swimtime="00:00:37.79"/><SPLIT distance="100" swimtime="00:01:21.41"/><SPLIT distance="150" swimtime="00:02:05.01"/></SPLITS></RESULT><RESULT eventid="10" heatid="150" lane="4" points="422" resultid="1133" swimtime="00:00:27.87"><SPLITS/></RESULT><RESULT eventid="12" heatid="184" lane="4" points="400" resultid="1392" swimtime="00:02:34.67"><SPLITS><SPLIT distance="50" swimtime="00:00:33.19"/><SPLIT distance="100" swimtime="00:01:15.58"/><SPLIT distance="150" swimtime="00:01:59.38"/></SPLITS></RESULT><RESULT eventid="32" heatid="354" lane="5" points="414" resultid="2639" swimtime="00:01:16.31"><SPLITS><SPLIT distance="50" swimtime="00:00:35.72"/></SPLITS></RESULT><RESULT eventid="40" heatid="470" lane="5" points="424" resultid="3518" swimtime="00:01:02.37"><SPLITS><SPLIT distance="50" swimtime="00:00:29.54"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="290" birthdate="2010-01-01" firstname="Pavel" gender="M" lastname="Gubanov" license="410664"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="38" lane="8" points="363" resultid="290" swimtime="00:00:36.35"><SPLITS/></RESULT><RESULT eventid="8" heatid="99" lane="4" points="354" resultid="744" swimtime="00:02:57.97"><SPLITS><SPLIT distance="50" swimtime="00:00:38.63"/><SPLIT distance="100" swimtime="00:01:24.40"/><SPLIT distance="150" swimtime="00:02:11.44"/></SPLITS></RESULT><RESULT eventid="10" heatid="147" lane="6" points="328" resultid="1111" swimtime="00:00:30.29"><SPLITS/></RESULT><RESULT eventid="12" heatid="184" lane="6" points="318" resultid="1393" swimtime="00:02:46.85"><SPLITS><SPLIT distance="50" swimtime="00:00:37.47"/><SPLIT distance="100" swimtime="00:01:22.90"/><SPLIT distance="150" swimtime="00:02:08.71"/></SPLITS></RESULT><RESULT eventid="28" heatid="282" lane="1" points="276" resultid="2093" swimtime="00:00:36.41"><SPLITS/></RESULT><RESULT eventid="32" heatid="354" lane="8" points="370" resultid="2642" swimtime="00:01:19.22"><SPLITS><SPLIT distance="50" swimtime="00:00:37.42"/></SPLITS></RESULT><RESULT eventid="36" heatid="391" lane="3" points="277" resultid="2912" swimtime="00:00:34.15"><SPLITS/></RESULT><RESULT eventid="40" heatid="466" lane="5" points="325" resultid="3487" swimtime="00:01:08.14"><SPLITS><SPLIT distance="50" swimtime="00:00:32.74"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="295" birthdate="2009-01-01" firstname="Lucas" gender="M" lastname="Platzer" license="416108"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="39" lane="5" points="526" resultid="295" swimtime="00:00:32.14"><SPLITS/></RESULT><RESULT eventid="8" heatid="100" lane="3" points="435" resultid="751" swimtime="00:02:46.10"><SPLITS><SPLIT distance="50" swimtime="00:00:37.11"/><SPLIT distance="100" swimtime="00:01:19.40"/><SPLIT distance="150" swimtime="00:02:04.07"/></SPLITS></RESULT><RESULT eventid="10" heatid="151" lane="2" points="408" resultid="1139" swimtime="00:00:28.17"><SPLITS/></RESULT><RESULT eventid="28" heatid="285" lane="7" points="388" resultid="2122" swimtime="00:00:32.49"><SPLITS/></RESULT><RESULT eventid="32" heatid="355" lane="2" points="471" resultid="2643" swimtime="00:01:13.07"><SPLITS><SPLIT distance="50" swimtime="00:00:33.66"/></SPLITS></RESULT><RESULT eventid="36" heatid="395" lane="6" points="396" resultid="2947" swimtime="00:00:30.32"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="298" birthdate="1998-01-01" firstname="Paul" gender="M" lastname="Deuker" license="248532"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="39" lane="8" points="346" resultid="298" swimtime="00:00:36.95"><SPLITS/></RESULT><RESULT eventid="10" heatid="156" lane="5" points="513" resultid="1180" swimtime="00:00:26.11"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="331" birthdate="2011-01-01" firstname="Mia" gender="F" lastname="Sibbe" license="495190"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="45" lane="4" points="253" resultid="339" swimtime="00:06:13.45"><SPLITS><SPLIT distance="100" swimtime="00:01:23.34"/><SPLIT distance="200" swimtime="00:02:59.09"/><SPLIT distance="300" swimtime="00:04:36.91"/></SPLITS></RESULT><RESULT eventid="9" heatid="118" lane="4" points="329" resultid="891" swimtime="00:00:34.27"><SPLITS/></RESULT><RESULT eventid="13" heatid="199" lane="5" points="220" resultid="1508" swimtime="00:01:35.13"><SPLITS><SPLIT distance="50" swimtime="00:00:44.39"/></SPLITS></RESULT><RESULT eventid="27" heatid="263" lane="8" points="184" resultid="1955" swimtime="00:00:47.42"><SPLITS/></RESULT><RESULT eventid="29" heatid="299" lane="3" points="262" resultid="2224" swimtime="00:02:56.53"><SPLITS><SPLIT distance="50" swimtime="00:00:38.71"/><SPLIT distance="100" swimtime="00:01:22.46"/><SPLIT distance="150" swimtime="00:02:11.13"/></SPLITS></RESULT><RESULT eventid="39" heatid="437" lane="5" resultid="3262" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="335" birthdate="2013-01-01" firstname="Emilia" gender="F" lastname="Paleani" license="451235"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="45" lane="8" points="323" resultid="343" swimtime="00:05:44.44"><SPLITS><SPLIT distance="100" swimtime="00:01:21.19"/><SPLIT distance="200" swimtime="00:02:48.81"/><SPLIT distance="300" swimtime="00:04:17.16"/></SPLITS></RESULT><RESULT eventid="9" heatid="115" lane="8" points="320" resultid="872" swimtime="00:00:34.58"><SPLITS/></RESULT><RESULT eventid="11" heatid="164" lane="6" points="334" resultid="1240" swimtime="00:03:01.68"><SPLITS><SPLIT distance="50" swimtime="00:00:38.00"/><SPLIT distance="100" swimtime="00:01:26.14"/><SPLIT distance="150" swimtime="00:02:21.50"/></SPLITS></RESULT><RESULT eventid="21" heatid="237" lane="4" resultid="1777" swimtime="00:00:55.21"><SPLITS/></RESULT><RESULT eventid="33" heatid="358" lane="2" points="267" resultid="2662" swimtime="00:03:09.08"><SPLITS><SPLIT distance="50" swimtime="00:00:41.19"/><SPLIT distance="100" swimtime="00:01:29.73"/><SPLIT distance="150" swimtime="00:02:20.66"/></SPLITS></RESULT><RESULT eventid="39" heatid="436" lane="7" points="325" resultid="3256" swimtime="00:01:15.15"><SPLITS><SPLIT distance="50" swimtime="00:00:36.48"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="363" birthdate="2009-01-01" firstname="Annika Lena" gender="F" lastname="Schwarz" license="416111"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="50" lane="8" points="435" resultid="382" swimtime="00:05:11.83"><SPLITS><SPLIT distance="100" swimtime="00:01:12.41"/><SPLIT distance="200" swimtime="00:02:32.76"/><SPLIT distance="300" swimtime="00:03:52.69"/></SPLITS></RESULT><RESULT eventid="9" heatid="128" lane="8" points="455" resultid="974" swimtime="00:00:30.77"><SPLITS/></RESULT><RESULT eventid="13" heatid="208" lane="7" points="450" resultid="1581" swimtime="00:01:14.94"><SPLITS><SPLIT distance="50" swimtime="00:00:36.13"/></SPLITS></RESULT><RESULT eventid="27" heatid="271" lane="1" points="457" resultid="2011" swimtime="00:00:35.02"><SPLITS/></RESULT><RESULT eventid="37" heatid="410" lane="2" points="448" resultid="3056" swimtime="00:02:41.18"><SPLITS><SPLIT distance="50" swimtime="00:00:37.28"/><SPLIT distance="100" swimtime="00:01:17.59"/><SPLIT distance="150" swimtime="00:01:59.91"/></SPLITS></RESULT><RESULT eventid="39" heatid="447" lane="3" points="483" resultid="3338" swimtime="00:01:05.87"><SPLITS><SPLIT distance="50" swimtime="00:00:32.08"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="368" birthdate="2008-01-01" firstname="Anna Maria" gender="F" lastname="Biernat" license="414127"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="51" lane="6" points="479" resultid="387" swimtime="00:05:01.98"><SPLITS><SPLIT distance="100" swimtime="00:01:10.88"/><SPLIT distance="200" swimtime="00:02:28.31"/><SPLIT distance="300" swimtime="00:03:46.16"/></SPLITS></RESULT><RESULT eventid="5" heatid="70" lane="1" points="428" resultid="520" swimtime="00:01:13.60"><SPLITS><SPLIT distance="50" swimtime="00:00:35.11"/></SPLITS></RESULT><RESULT eventid="9" heatid="128" lane="2" points="478" resultid="968" swimtime="00:00:30.27"><SPLITS/></RESULT><RESULT eventid="11" heatid="172" lane="4" points="487" resultid="1302" swimtime="00:02:40.30"><SPLITS><SPLIT distance="50" swimtime="00:00:32.57"/><SPLIT distance="100" swimtime="00:01:16.47"/><SPLIT distance="150" swimtime="00:02:03.62"/></SPLITS></RESULT><RESULT eventid="29" heatid="306" lane="1" points="481" resultid="2275" swimtime="00:02:24.19"><SPLITS><SPLIT distance="50" swimtime="00:00:32.58"/><SPLIT distance="100" swimtime="00:01:08.48"/><SPLIT distance="150" swimtime="00:01:46.42"/></SPLITS></RESULT><RESULT eventid="35" heatid="380" lane="2" resultid="2829" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="39" heatid="448" lane="8" resultid="3350" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="372" birthdate="2010-01-01" firstname="Noemi" gender="F" lastname="Varga" license="422346"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="52" lane="2" points="486" resultid="391" swimtime="00:05:00.61"><SPLITS><SPLIT distance="100" swimtime="00:01:08.78"/><SPLIT distance="200" swimtime="00:02:24.60"/><SPLIT distance="300" swimtime="00:03:42.79"/></SPLITS></RESULT><RESULT comment="15:54 Die Sportlerin hat beim Abstoß bei der Teilstrecke Brust die Bahn verlassen" eventid="11" heatid="171" lane="6" resultid="1296" status="DSQ" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="17" heatid="231" lane="4" points="495" resultid="1743" swimtime="00:10:12.67"><SPLITS><SPLIT distance="100" swimtime="00:01:09.03"/><SPLIT distance="200" swimtime="00:02:24.23"/><SPLIT distance="300" swimtime="00:03:40.58"/><SPLIT distance="400" swimtime="00:04:58.73"/><SPLIT distance="500" swimtime="00:06:16.91"/><SPLIT distance="600" swimtime="00:07:35.90"/><SPLIT distance="700" swimtime="00:08:55.00"/></SPLITS></RESULT><RESULT eventid="29" heatid="306" lane="5" points="475" resultid="2279" swimtime="00:02:24.78"><SPLITS><SPLIT distance="50" swimtime="00:00:33.08"/><SPLIT distance="100" swimtime="00:01:09.45"/><SPLIT distance="150" swimtime="00:01:47.21"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="395" birthdate="2015-01-01" firstname="Benedikt" gender="M" lastname="Maierhofer" license="454097"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="56" lane="2" points="182" resultid="419" swimtime="00:06:27.98"><SPLITS><SPLIT distance="100" swimtime="00:01:29.53"/><SPLIT distance="200" swimtime="00:03:12.06"/><SPLIT distance="300" swimtime="00:04:52.85"/></SPLITS></RESULT><RESULT eventid="10" heatid="144" lane="1" points="170" resultid="1082" swimtime="00:00:37.68"><SPLITS/></RESULT><RESULT eventid="14" heatid="217" lane="7" points="153" resultid="1649" swimtime="00:01:36.44"><SPLITS><SPLIT distance="50" swimtime="00:00:47.19"/></SPLITS></RESULT><RESULT eventid="30" heatid="315" lane="5" points="162" resultid="2346" swimtime="00:03:06.92"><SPLITS><SPLIT distance="50" swimtime="00:00:40.05"/><SPLIT distance="100" swimtime="00:01:29.63"/><SPLIT distance="150" swimtime="00:02:19.38"/></SPLITS></RESULT><RESULT eventid="32" heatid="347" lane="2" points="106" resultid="2583" swimtime="00:02:00.00"><SPLITS><SPLIT distance="50" swimtime="00:00:57.35"/></SPLITS></RESULT><RESULT eventid="36" heatid="386" lane="6" points="88" resultid="2876" swimtime="00:00:49.93"><SPLITS/></RESULT><RESULT eventid="40" heatid="460" lane="5" points="154" resultid="3440" swimtime="00:01:27.39"><SPLITS><SPLIT distance="50" swimtime="00:00:41.80"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="406" birthdate="2014-01-01" firstname="Jasim" gender="M" lastname="Al-Sultan" license="449445"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="57" lane="8" points="234" resultid="433" swimtime="00:05:56.79"><SPLITS><SPLIT distance="100" swimtime="00:01:23.94"/><SPLIT distance="200" swimtime="00:02:56.00"/><SPLIT distance="300" swimtime="00:04:28.15"/></SPLITS></RESULT><RESULT eventid="8" heatid="93" lane="5" points="152" resultid="701" swimtime="00:03:55.81"><SPLITS><SPLIT distance="50" swimtime="00:00:54.13"/><SPLIT distance="100" swimtime="00:01:55.82"/><SPLIT distance="150" swimtime="00:02:55.52"/></SPLITS></RESULT><RESULT eventid="12" heatid="177" lane="8" points="166" resultid="1342" swimtime="00:03:27.30"><SPLITS><SPLIT distance="50" swimtime="00:00:57.18"/><SPLIT distance="100" swimtime="00:01:45.38"/><SPLIT distance="150" swimtime="00:02:44.57"/></SPLITS></RESULT><RESULT eventid="24" heatid="244" lane="2" resultid="1815" swimtime="00:00:58.33"><SPLITS/></RESULT><RESULT eventid="30" heatid="316" lane="1" points="206" resultid="2350" swimtime="00:02:52.62"><SPLITS><SPLIT distance="50" swimtime="00:00:40.24"/><SPLIT distance="100" swimtime="00:01:24.41"/><SPLIT distance="150" swimtime="00:02:09.82"/></SPLITS></RESULT><RESULT eventid="32" heatid="347" lane="7" points="116" resultid="2588" swimtime="00:01:56.55"><SPLITS><SPLIT distance="50" swimtime="00:00:55.78"/></SPLITS></RESULT><RESULT eventid="40" heatid="459" lane="5" points="176" resultid="3433" swimtime="00:01:23.54"><SPLITS><SPLIT distance="50" swimtime="00:00:39.62"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="408" birthdate="2013-01-01" firstname="Levin" gender="M" lastname="Burkhart" license="452028"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="58" lane="3" points="253" resultid="436" swimtime="00:05:47.50"><SPLITS><SPLIT distance="100" swimtime="00:01:19.68"/><SPLIT distance="200" swimtime="00:02:50.08"/><SPLIT distance="300" swimtime="00:04:20.86"/></SPLITS></RESULT><RESULT eventid="12" heatid="180" lane="8" points="224" resultid="1365" swimtime="00:03:07.48"><SPLITS><SPLIT distance="50" swimtime="00:00:45.78"/><SPLIT distance="100" swimtime="00:01:30.58"/><SPLIT distance="150" swimtime="00:02:29.14"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="413" birthdate="2013-01-01" firstname="Viktor" gender="M" lastname="Gubanov" license="422857"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="59" lane="2" points="348" resultid="442" swimtime="00:05:12.79"><SPLITS><SPLIT distance="100" swimtime="00:01:12.79"/><SPLIT distance="200" swimtime="00:02:32.90"/><SPLIT distance="300" swimtime="00:03:54.50"/></SPLITS></RESULT><RESULT eventid="12" heatid="183" lane="4" points="300" resultid="1385" swimtime="00:02:50.27"><SPLITS><SPLIT distance="50" swimtime="00:00:35.68"/><SPLIT distance="100" swimtime="00:01:21.50"/><SPLIT distance="150" swimtime="00:02:12.77"/></SPLITS></RESULT><RESULT eventid="20" heatid="236" lane="6" resultid="1774" swimtime="00:00:46.00"><SPLITS/></RESULT><RESULT eventid="30" heatid="320" lane="7" points="327" resultid="2388" swimtime="00:02:27.95"><SPLITS><SPLIT distance="50" swimtime="00:00:33.19"/><SPLIT distance="100" swimtime="00:01:11.56"/><SPLIT distance="150" swimtime="00:01:50.56"/></SPLITS></RESULT><RESULT eventid="38" heatid="418" lane="8" points="264" resultid="3120" swimtime="00:02:54.30"><SPLITS><SPLIT distance="50" swimtime="00:00:40.55"/><SPLIT distance="100" swimtime="00:01:25.06"/><SPLIT distance="150" swimtime="00:02:10.68"/></SPLITS></RESULT><RESULT eventid="40" heatid="467" lane="7" points="305" resultid="3496" swimtime="00:01:09.58"><SPLITS><SPLIT distance="50" swimtime="00:00:32.07"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="423" birthdate="2011-01-01" firstname="Niklas" gender="M" lastname="Luber" license="407350"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="60" lane="4" points="424" resultid="452" swimtime="00:04:52.85"><SPLITS><SPLIT distance="100" swimtime="00:01:07.87"/><SPLIT distance="200" swimtime="00:02:22.65"/><SPLIT distance="300" swimtime="00:03:37.89"/></SPLITS></RESULT><RESULT eventid="18" heatid="233" lane="8" points="413" resultid="1758" swimtime="00:10:06.92"><SPLITS><SPLIT distance="100" swimtime="00:01:07.57"/><SPLIT distance="200" swimtime="00:02:23.66"/><SPLIT distance="300" swimtime="00:03:41.31"/><SPLIT distance="400" swimtime="00:04:57.89"/><SPLIT distance="500" swimtime="00:06:15.88"/><SPLIT distance="600" swimtime="00:07:33.81"/><SPLIT distance="700" swimtime="00:08:50.78"/></SPLITS></RESULT><RESULT eventid="30" heatid="323" lane="1" points="403" resultid="2404" swimtime="00:02:18.03"><SPLITS><SPLIT distance="50" swimtime="00:00:30.67"/><SPLIT distance="100" swimtime="00:01:05.27"/><SPLIT distance="150" swimtime="00:01:42.24"/></SPLITS></RESULT><RESULT eventid="40" heatid="470" lane="1" points="406" resultid="3514" swimtime="00:01:03.27"><SPLITS><SPLIT distance="50" swimtime="00:00:30.83"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="430" birthdate="2010-01-01" firstname="Maxim" gender="M" lastname="Frenkel" license="397963"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="61" lane="4" points="497" resultid="459" swimtime="00:04:37.75"><SPLITS><SPLIT distance="100" swimtime="00:01:02.93"/><SPLIT distance="200" swimtime="00:02:13.78"/><SPLIT distance="300" swimtime="00:03:26.53"/></SPLITS></RESULT><RESULT eventid="10" heatid="150" lane="2" points="422" resultid="1131" swimtime="00:00:27.87"><SPLITS/></RESULT><RESULT eventid="12" heatid="189" lane="1" points="482" resultid="1428" swimtime="00:02:25.34"><SPLITS><SPLIT distance="50" swimtime="00:00:31.62"/><SPLIT distance="100" swimtime="00:01:08.97"/><SPLIT distance="150" swimtime="00:01:52.11"/></SPLITS></RESULT><RESULT eventid="30" heatid="324" lane="1" points="493" resultid="2411" swimtime="00:02:09.11"><SPLITS><SPLIT distance="50" swimtime="00:00:29.77"/><SPLIT distance="100" swimtime="00:01:02.03"/><SPLIT distance="150" swimtime="00:01:36.07"/></SPLITS></RESULT><RESULT eventid="40" heatid="470" lane="7" points="477" resultid="3520" swimtime="00:00:59.96"><SPLITS><SPLIT distance="50" swimtime="00:00:28.54"/></SPLITS></RESULT><RESULT eventid="42" heatid="481" lane="7" points="477" resultid="3596" swimtime="00:05:12.01"><SPLITS><SPLIT distance="50" swimtime="00:00:32.21"/><SPLIT distance="100" swimtime="00:01:11.55"/><SPLIT distance="150" swimtime="00:01:50.05"/><SPLIT distance="200" swimtime="00:02:30.00"/><SPLIT distance="250" swimtime="00:03:15.69"/><SPLIT distance="300" swimtime="00:04:01.74"/><SPLIT distance="350" swimtime="00:04:37.26"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="437" birthdate="2009-01-01" firstname="Julius" gender="M" lastname="Tokaji" license="436951"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="62" lane="7" points="539" resultid="467" swimtime="00:04:30.27"><SPLITS><SPLIT distance="100" swimtime="00:01:03.92"/><SPLIT distance="200" swimtime="00:02:13.06"/><SPLIT distance="300" swimtime="00:03:22.31"/></SPLITS></RESULT><RESULT eventid="18" heatid="233" lane="4" points="529" resultid="1755" swimtime="00:09:18.88"><SPLITS><SPLIT distance="100" swimtime="00:01:04.69"/><SPLIT distance="200" swimtime="00:02:14.69"/><SPLIT distance="300" swimtime="00:03:25.07"/><SPLIT distance="400" swimtime="00:04:35.83"/><SPLIT distance="500" swimtime="00:05:46.83"/><SPLIT distance="600" swimtime="00:06:57.80"/><SPLIT distance="700" swimtime="00:08:09.05"/></SPLITS></RESULT><RESULT eventid="30" heatid="324" lane="8" points="532" resultid="2418" swimtime="00:02:05.88"><SPLITS><SPLIT distance="50" swimtime="00:00:29.66"/><SPLIT distance="100" swimtime="00:01:00.88"/><SPLIT distance="150" swimtime="00:01:34.12"/></SPLITS></RESULT><RESULT eventid="40" heatid="471" lane="5" points="529" resultid="3526" swimtime="00:00:57.91"><SPLITS><SPLIT distance="50" swimtime="00:00:28.10"/></SPLITS></RESULT><RESULT eventid="42" heatid="479" lane="2" points="468" resultid="3579" swimtime="00:05:14.00"><SPLITS><SPLIT distance="50" swimtime="00:00:32.48"/><SPLIT distance="100" swimtime="00:01:11.06"/><SPLIT distance="150" swimtime="00:01:53.10"/><SPLIT distance="200" swimtime="00:02:33.00"/><SPLIT distance="250" swimtime="00:03:18.54"/><SPLIT distance="300" swimtime="00:04:03.74"/><SPLIT distance="350" swimtime="00:04:39.80"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="445" birthdate="2013-01-01" firstname="Lisa" gender="F" lastname="Weizel" license="436957"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="5" heatid="65" lane="4" points="237" resultid="484" swimtime="00:01:29.65"><SPLITS><SPLIT distance="50" swimtime="00:00:39.69"/></SPLITS></RESULT><RESULT eventid="11" heatid="167" lane="8" points="332" resultid="1266" swimtime="00:03:02.04"><SPLITS><SPLIT distance="50" swimtime="00:00:41.80"/><SPLIT distance="100" swimtime="00:01:26.49"/><SPLIT distance="150" swimtime="00:02:21.53"/></SPLITS></RESULT><RESULT eventid="13" heatid="201" lane="1" points="312" resultid="1520" swimtime="00:01:24.69"><SPLITS><SPLIT distance="50" swimtime="00:00:42.26"/></SPLITS></RESULT><RESULT eventid="21" heatid="237" lane="5" resultid="1778" swimtime="00:00:57.13"><SPLITS/></RESULT><RESULT eventid="39" heatid="436" lane="3" points="312" resultid="3252" swimtime="00:01:16.22"><SPLITS><SPLIT distance="50" swimtime="00:00:36.30"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="457" birthdate="2009-01-01" firstname="Martha" gender="F" lastname="Albrecht" license="380190"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="5" heatid="69" lane="4" points="496" resultid="515" swimtime="00:01:10.07"><SPLITS><SPLIT distance="50" swimtime="00:00:30.60"/></SPLITS></RESULT><RESULT eventid="7" heatid="92" lane="8" points="527" resultid="696" swimtime="00:02:52.00"><SPLITS><SPLIT distance="50" swimtime="00:00:39.13"/><SPLIT distance="100" swimtime="00:01:22.47"/><SPLIT distance="150" swimtime="00:02:08.36"/></SPLITS></RESULT><RESULT eventid="11" heatid="172" lane="6" points="495" resultid="1304" swimtime="00:02:39.40"><SPLITS><SPLIT distance="50" swimtime="00:00:32.22"/><SPLIT distance="100" swimtime="00:01:14.77"/><SPLIT distance="150" swimtime="00:02:00.59"/></SPLITS></RESULT><RESULT eventid="31" heatid="344" lane="1" points="559" resultid="2563" swimtime="00:01:17.84"><SPLITS><SPLIT distance="50" swimtime="00:00:37.80"/></SPLITS></RESULT><RESULT eventid="35" heatid="382" lane="1" points="519" resultid="2844" swimtime="00:00:30.39"><SPLITS/></RESULT><RESULT eventid="37" heatid="410" lane="7" points="448" resultid="3061" swimtime="00:02:41.12"><SPLITS><SPLIT distance="50" swimtime="00:00:36.76"/><SPLIT distance="100" swimtime="00:01:17.89"/><SPLIT distance="150" swimtime="00:01:59.69"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="458" birthdate="2011-01-01" firstname="Sophie" gender="F" lastname="Nibler" license="421036"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="5" heatid="69" lane="7" resultid="518" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="9" heatid="124" lane="2" resultid="937" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="11" heatid="168" lane="1" resultid="1267" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="27" heatid="267" lane="8" points="290" resultid="1987" swimtime="00:00:40.72"><SPLITS/></RESULT><RESULT eventid="29" heatid="301" lane="6" points="413" resultid="2242" swimtime="00:02:31.62"><SPLITS><SPLIT distance="50" swimtime="00:00:34.66"/><SPLIT distance="100" swimtime="00:01:12.78"/><SPLIT distance="150" swimtime="00:01:52.92"/></SPLITS></RESULT><RESULT eventid="33" heatid="358" lane="3" points="308" resultid="2663" swimtime="00:03:00.24"><SPLITS><SPLIT distance="50" swimtime="00:00:36.44"/><SPLIT distance="100" swimtime="00:01:20.81"/><SPLIT distance="150" swimtime="00:02:10.07"/></SPLITS></RESULT><RESULT eventid="35" heatid="378" lane="4" points="397" resultid="2815" swimtime="00:00:33.22"><SPLITS/></RESULT><RESULT eventid="39" heatid="442" lane="6" points="405" resultid="3302" swimtime="00:01:09.89"><SPLITS><SPLIT distance="50" swimtime="00:00:33.91"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="495" birthdate="2009-01-01" firstname="Oliver" gender="M" lastname="Priese" license="422363"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="6" heatid="78" lane="5" points="471" resultid="586" swimtime="00:01:03.53"><SPLITS><SPLIT distance="50" swimtime="00:00:28.93"/></SPLITS></RESULT><RESULT eventid="10" heatid="155" lane="7" points="530" resultid="1174" swimtime="00:00:25.83"><SPLITS/></RESULT><RESULT eventid="36" heatid="399" lane="1" points="521" resultid="2974" swimtime="00:00:27.67"><SPLITS/></RESULT><RESULT eventid="40" heatid="473" lane="5" points="560" resultid="3541" swimtime="00:00:56.83"><SPLITS><SPLIT distance="50" swimtime="00:00:27.52"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="496" birthdate="2009-01-01" firstname="Jakub" gender="M" lastname="Vitkovic" license="422343"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="6" heatid="78" lane="8" points="412" resultid="589" swimtime="00:01:06.41"><SPLITS><SPLIT distance="50" swimtime="00:00:30.63"/></SPLITS></RESULT><RESULT eventid="10" heatid="151" lane="5" points="448" resultid="1142" swimtime="00:00:27.32"><SPLITS/></RESULT><RESULT eventid="14" heatid="224" lane="2" points="443" resultid="1698" swimtime="00:01:07.65"><SPLITS><SPLIT distance="50" swimtime="00:00:32.73"/></SPLITS></RESULT><RESULT comment="09:47 Start vor dem Startsignal" eventid="28" heatid="286" lane="1" resultid="2124" status="DSQ" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="30" heatid="323" lane="7" points="505" resultid="2409" swimtime="00:02:08.07"><SPLITS><SPLIT distance="50" swimtime="00:00:28.75"/><SPLIT distance="100" swimtime="00:01:01.88"/><SPLIT distance="150" swimtime="00:01:35.80"/></SPLITS></RESULT><RESULT eventid="36" heatid="397" lane="8" points="424" resultid="2965" swimtime="00:00:29.63"><SPLITS/></RESULT><RESULT eventid="40" heatid="471" lane="3" points="534" resultid="3524" swimtime="00:00:57.74"><SPLITS><SPLIT distance="50" swimtime="00:00:28.16"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="506" birthdate="2013-01-01" firstname="Anna" gender="F" lastname="Weizel" license="436958"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="7" heatid="87" lane="3" points="343" resultid="651" swimtime="00:03:18.31"><SPLITS><SPLIT distance="50" swimtime="00:00:44.77"/><SPLIT distance="100" swimtime="00:01:35.96"/><SPLIT distance="150" swimtime="00:02:27.87"/></SPLITS></RESULT><RESULT eventid="11" heatid="167" lane="7" points="357" resultid="1265" swimtime="00:02:57.71"><SPLITS><SPLIT distance="50" swimtime="00:00:41.98"/><SPLIT distance="100" swimtime="00:01:27.95"/><SPLIT distance="150" swimtime="00:02:17.82"/></SPLITS></RESULT><RESULT eventid="25" heatid="247" lane="6" resultid="1835" swimtime="00:00:59.24"><SPLITS/></RESULT><RESULT eventid="31" heatid="339" lane="8" points="332" resultid="2530" swimtime="00:01:32.54"><SPLITS><SPLIT distance="50" swimtime="00:00:44.39"/></SPLITS></RESULT><RESULT eventid="37" heatid="406" lane="2" points="330" resultid="3024" swimtime="00:02:58.32"><SPLITS><SPLIT distance="50" swimtime="00:00:42.85"/><SPLIT distance="100" swimtime="00:01:27.43"/><SPLIT distance="150" swimtime="00:02:14.09"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="511" birthdate="2015-01-01" firstname="Elias" gender="M" lastname="Henkel" license="461538"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="8" heatid="95" lane="7" points="173" resultid="716" swimtime="00:03:45.66"><SPLITS><SPLIT distance="50" swimtime="00:00:51.76"/><SPLIT distance="100" swimtime="00:01:50.18"/><SPLIT distance="150" swimtime="00:02:49.79"/></SPLITS></RESULT><RESULT eventid="10" heatid="141" lane="1" points="125" resultid="1059" swimtime="00:00:41.82"><SPLITS/></RESULT><RESULT eventid="12" heatid="175" lane="3" points="146" resultid="1324" swimtime="00:03:36.09"><SPLITS><SPLIT distance="50" swimtime="00:00:54.79"/><SPLIT distance="100" swimtime="00:01:47.48"/><SPLIT distance="150" swimtime="00:02:45.66"/></SPLITS></RESULT><RESULT eventid="14" heatid="215" lane="3" points="123" resultid="1630" swimtime="00:01:43.75"><SPLITS><SPLIT distance="50" swimtime="00:00:52.14"/></SPLITS></RESULT><RESULT eventid="30" heatid="311" lane="5" points="142" resultid="2316" swimtime="00:03:15.22"><SPLITS><SPLIT distance="50" swimtime="00:00:43.37"/><SPLIT distance="100" swimtime="00:01:34.87"/><SPLIT distance="150" swimtime="00:02:26.71"/></SPLITS></RESULT><RESULT eventid="32" heatid="349" lane="2" points="147" resultid="2598" swimtime="00:01:47.74"><SPLITS><SPLIT distance="50" swimtime="00:00:51.25"/></SPLITS></RESULT><RESULT eventid="36" heatid="387" lane="7" points="91" resultid="2884" swimtime="00:00:49.41"><SPLITS/></RESULT><RESULT eventid="40" heatid="458" lane="1" points="135" resultid="3421" swimtime="00:01:31.30"><SPLITS><SPLIT distance="50" swimtime="00:00:42.88"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="513" birthdate="2015-01-01" firstname="Johanna" gender="F" lastname="Enneking" license="472022"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="9" heatid="106" lane="4" points="194" resultid="796" swimtime="00:00:40.83"><SPLITS/></RESULT><RESULT eventid="13" heatid="191" lane="8" points="136" resultid="1447" swimtime="00:01:51.51"><SPLITS><SPLIT distance="50" swimtime="00:00:54.09"/></SPLITS></RESULT><RESULT eventid="31" heatid="327" lane="4" points="150" resultid="2431" swimtime="00:02:00.65"><SPLITS><SPLIT distance="50" swimtime="00:00:56.56"/></SPLITS></RESULT><RESULT eventid="35" heatid="365" lane="6" points="114" resultid="2716" swimtime="00:00:50.37"><SPLITS/></RESULT><RESULT eventid="39" heatid="423" lane="7" points="126" resultid="3153" swimtime="00:01:42.96"><SPLITS><SPLIT distance="50" swimtime="00:00:45.90"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="522" birthdate="2005-01-01" firstname="Jana" gender="F" lastname="Said" license="416384"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="9" heatid="121" lane="1" points="364" resultid="912" swimtime="00:00:33.13"><SPLITS/></RESULT><RESULT eventid="13" heatid="205" lane="5" points="398" resultid="1556" swimtime="00:01:18.09"><SPLITS><SPLIT distance="50" swimtime="00:00:37.58"/></SPLITS></RESULT><RESULT eventid="27" heatid="269" lane="5" points="424" resultid="1999" swimtime="00:00:35.90"><SPLITS/></RESULT><RESULT eventid="37" heatid="408" lane="4" points="399" resultid="3042" swimtime="00:02:47.51"><SPLITS><SPLIT distance="50" swimtime="00:00:39.31"/><SPLIT distance="100" swimtime="00:01:22.47"/><SPLIT distance="150" swimtime="00:02:04.84"/></SPLITS></RESULT><RESULT eventid="39" heatid="439" lane="1" points="357" resultid="3274" swimtime="00:01:12.88"><SPLITS><SPLIT distance="50" swimtime="00:00:35.21"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="527" birthdate="2007-01-01" firstname="Eleonora" gender="F" lastname="van de Kuilen" license="432200"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="9" heatid="125" lane="2" points="456" resultid="945" swimtime="00:00:30.74"><SPLITS/></RESULT><RESULT eventid="13" heatid="202" lane="6" points="335" resultid="1533" swimtime="00:01:22.65"><SPLITS><SPLIT distance="50" swimtime="00:00:40.14"/></SPLITS></RESULT><RESULT eventid="27" heatid="265" lane="4" points="366" resultid="1967" swimtime="00:00:37.71"><SPLITS/></RESULT><RESULT eventid="29" heatid="301" lane="1" points="401" resultid="2238" swimtime="00:02:33.10"><SPLITS><SPLIT distance="50" swimtime="00:00:35.83"/><SPLIT distance="100" swimtime="00:01:13.98"/><SPLIT distance="150" swimtime="00:01:54.64"/></SPLITS></RESULT><RESULT eventid="35" heatid="373" lane="3" points="333" resultid="2777" swimtime="00:00:35.23"><SPLITS/></RESULT><RESULT eventid="39" heatid="443" lane="6" points="414" resultid="3310" swimtime="00:01:09.37"><SPLITS><SPLIT distance="50" swimtime="00:00:33.13"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="557" birthdate="2008-01-01" firstname="Max" gender="M" lastname="Rottmann" license="412987"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="10" heatid="154" lane="8" resultid="1168" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="14" heatid="224" lane="7" resultid="1703" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="28" heatid="286" lane="6" resultid="2129" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="36" heatid="397" lane="3" resultid="2960" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="559" birthdate="2003-01-01" firstname="Huba" gender="M" lastname="Pathi" license="303293"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="10" heatid="156" lane="4" resultid="1179" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="14" heatid="225" lane="3" resultid="1706" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="28" heatid="287" lane="3" points="504" resultid="2134" swimtime="00:00:29.79"><SPLITS/></RESULT><RESULT eventid="36" heatid="400" lane="6" points="498" resultid="2986" swimtime="00:00:28.08"><SPLITS/></RESULT><RESULT eventid="40" heatid="474" lane="6" points="523" resultid="3550" swimtime="00:00:58.15"><SPLITS><SPLIT distance="50" swimtime="00:00:27.45"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="568" birthdate="2002-01-01" firstname="Niklas" gender="M" lastname="Ludwig" license="486359"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="16" heatid="229" lane="3" points="562" resultid="1727" swimtime="00:17:35.01"><SPLITS><SPLIT distance="100" swimtime="00:01:05.40"/><SPLIT distance="200" swimtime="00:02:15.56"/><SPLIT distance="300" swimtime="00:03:26.22"/><SPLIT distance="400" swimtime="00:04:37.14"/><SPLIT distance="500" swimtime="00:05:48.23"/><SPLIT distance="600" swimtime="00:06:58.99"/><SPLIT distance="700" swimtime="00:08:10.01"/><SPLIT distance="800" swimtime="00:09:20.85"/><SPLIT distance="900" swimtime="00:10:31.74"/><SPLIT distance="1000" swimtime="00:11:42.73"/><SPLIT distance="1100" swimtime="00:12:53.48"/><SPLIT distance="1200" swimtime="00:14:04.05"/><SPLIT distance="1300" swimtime="00:15:15.18"/><SPLIT distance="1400" swimtime="00:16:26.18"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="578" birthdate="2013-01-01" firstname="Katharina" gender="F" lastname="Schmidt" license="497256"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="27" heatid="260" lane="1" points="200" resultid="1924" swimtime="00:00:46.09"><SPLITS/></RESULT><RESULT eventid="29" heatid="291" lane="7" points="193" resultid="2164" swimtime="00:03:15.33"><SPLITS><SPLIT distance="50" swimtime="00:00:41.70"/><SPLIT distance="100" swimtime="00:01:33.71"/><SPLIT distance="150" swimtime="00:02:26.55"/></SPLITS></RESULT><RESULT eventid="37" heatid="402" lane="4" points="184" resultid="2995" swimtime="00:03:36.73"><SPLITS><SPLIT distance="50" swimtime="00:00:49.21"/><SPLIT distance="100" swimtime="00:01:47.09"/><SPLIT distance="150" swimtime="00:02:43.44"/></SPLITS></RESULT><RESULT eventid="39" heatid="424" lane="1" points="171" resultid="3155" swimtime="00:01:33.14"><SPLITS><SPLIT distance="50" swimtime="00:00:45.42"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="579" birthdate="2015-01-01" firstname="Paula" gender="F" lastname="Seiwert" license="470828"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="27" heatid="260" lane="2" points="199" resultid="1925" swimtime="00:00:46.19"><SPLITS/></RESULT><RESULT eventid="29" heatid="293" lane="3" points="241" resultid="2176" swimtime="00:03:01.48"><SPLITS><SPLIT distance="50" swimtime="00:00:42.18"/><SPLIT distance="100" swimtime="00:01:27.96"/><SPLIT distance="150" swimtime="00:02:15.74"/></SPLITS></RESULT><RESULT eventid="31" heatid="332" lane="2" points="174" resultid="2468" swimtime="00:01:54.87"><SPLITS><SPLIT distance="50" swimtime="00:00:55.98"/></SPLITS></RESULT><RESULT eventid="35" heatid="367" lane="8" points="131" resultid="2734" swimtime="00:00:48.05"><SPLITS/></RESULT><RESULT eventid="39" heatid="426" lane="5" points="222" resultid="3174" swimtime="00:01:25.31"><SPLITS><SPLIT distance="50" swimtime="00:00:39.21"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="581" birthdate="2012-01-01" firstname="Polina" gender="F" lastname="Zinkevych" license="460352"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="27" heatid="263" lane="4" points="273" resultid="1951" swimtime="00:00:41.55"><SPLITS/></RESULT><RESULT eventid="31" heatid="340" lane="5" points="322" resultid="2535" swimtime="00:01:33.49"><SPLITS><SPLIT distance="50" swimtime="00:00:44.33"/></SPLITS></RESULT><RESULT eventid="35" heatid="370" lane="4" points="231" resultid="2754" swimtime="00:00:39.76"><SPLITS/></RESULT><RESULT eventid="39" heatid="436" lane="5" points="297" resultid="3254" swimtime="00:01:17.45"><SPLITS><SPLIT distance="50" swimtime="00:00:37.05"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="587" birthdate="2009-01-01" firstname="Sarah" gender="F" lastname="Obieglo" license="359759"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="27" heatid="271" lane="4" resultid="2013" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="29" heatid="306" lane="3" resultid="2277" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="35" heatid="377" lane="6" resultid="2810" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="37" heatid="411" lane="5" resultid="3067" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="39" heatid="449" lane="1" resultid="3351" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="592" birthdate="2014-01-01" firstname="Gabriel" gender="M" lastname="Sannino Murakame" license="501517"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="28" heatid="276" lane="2" points="81" resultid="2048" swimtime="00:00:54.66"><SPLITS/></RESULT><RESULT comment="12:43 Der Sportler verließ nach der 50m Wende die Wand bevor er vollständig in die Bauchlage zurückgekehrt war" eventid="32" heatid="347" lane="8" resultid="2589" status="DSQ" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="40" heatid="455" lane="6" points="107" resultid="3403" swimtime="00:01:38.51"><SPLITS><SPLIT distance="50" swimtime="00:00:45.92"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="595" birthdate="2015-01-01" firstname="Quentin" gender="M" lastname="Domurado" license="467535"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="28" heatid="280" lane="8" points="136" resultid="2084" swimtime="00:00:46.08"><SPLITS/></RESULT><RESULT eventid="30" heatid="314" lane="1" points="184" resultid="2334" swimtime="00:02:59.06"><SPLITS><SPLIT distance="50" swimtime="00:00:40.59"/><SPLIT distance="100" swimtime="00:01:28.62"/><SPLIT distance="150" swimtime="00:02:15.06"/></SPLITS></RESULT><RESULT eventid="32" heatid="348" lane="4" points="127" resultid="2593" swimtime="00:01:52.91"><SPLITS><SPLIT distance="50" swimtime="00:00:53.49"/></SPLITS></RESULT><RESULT eventid="36" heatid="388" lane="5" points="123" resultid="2890" swimtime="00:00:44.68"><SPLITS/></RESULT><RESULT eventid="38" heatid="415" lane="6" points="170" resultid="3096" swimtime="00:03:22.02"><SPLITS><SPLIT distance="50" swimtime="00:00:48.38"/><SPLIT distance="100" swimtime="00:01:40.53"/><SPLIT distance="150" swimtime="00:02:32.61"/></SPLITS></RESULT><RESULT eventid="40" heatid="459" lane="2" points="146" resultid="3430" swimtime="00:01:28.87"><SPLITS><SPLIT distance="50" swimtime="00:00:43.24"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="598" birthdate="2010-01-01" firstname="Jonas" gender="M" lastname="Scheffel" license="435049"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="28" heatid="287" lane="8" points="437" resultid="2137" swimtime="00:00:31.24"><SPLITS/></RESULT><RESULT eventid="36" heatid="398" lane="4" points="508" resultid="2969" swimtime="00:00:27.90"><SPLITS/></RESULT><RESULT eventid="40" heatid="473" lane="6" points="495" resultid="3542" swimtime="00:00:59.20"><SPLITS><SPLIT distance="50" swimtime="00:00:28.81"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="599" birthdate="2012-01-01" firstname="Magdalena" gender="F" lastname="Bär" license="436952"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="29" heatid="303" lane="4" points="516" resultid="2256" swimtime="00:02:20.81"><SPLITS><SPLIT distance="50" swimtime="00:00:33.08"/><SPLIT distance="100" swimtime="00:01:09.08"/><SPLIT distance="150" swimtime="00:01:45.13"/></SPLITS></RESULT><RESULT eventid="35" heatid="376" lane="1" points="403" resultid="2798" swimtime="00:00:33.06"><SPLITS/></RESULT><RESULT eventid="37" heatid="411" lane="8" points="470" resultid="3070" swimtime="00:02:38.63"><SPLITS><SPLIT distance="100" swimtime="00:01:17.23"/></SPLITS></RESULT><RESULT eventid="39" heatid="445" lane="5" points="481" resultid="3325" swimtime="00:01:05.98"><SPLITS><SPLIT distance="50" swimtime="00:00:32.22"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="600" birthdate="2006-01-01" firstname="Johanna Marie" gender="F" lastname="Schwarz" license="416112"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="29" heatid="304" lane="5" points="384" resultid="2265" swimtime="00:02:35.37"><SPLITS><SPLIT distance="50" swimtime="00:00:34.53"/><SPLIT distance="100" swimtime="00:01:13.09"/><SPLIT distance="150" swimtime="00:01:55.26"/></SPLITS></RESULT><RESULT eventid="39" heatid="446" lane="3" points="400" resultid="3330" swimtime="00:01:10.17"><SPLITS><SPLIT distance="50" swimtime="00:00:33.84"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="601" birthdate="2008-01-01" firstname="Maria" gender="F" lastname="Obieglo" license="351446"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="29" heatid="307" lane="1" points="532" resultid="2283" swimtime="00:02:19.37"><SPLITS><SPLIT distance="50" swimtime="00:00:33.45"/><SPLIT distance="100" swimtime="00:01:08.30"/><SPLIT distance="150" swimtime="00:01:44.99"/></SPLITS></RESULT><RESULT eventid="33" heatid="360" lane="5" points="488" resultid="2679" swimtime="00:02:34.68"><SPLITS><SPLIT distance="50" swimtime="00:00:34.33"/><SPLIT distance="100" swimtime="00:01:12.60"/><SPLIT distance="150" swimtime="00:01:53.35"/></SPLITS></RESULT><RESULT eventid="35" heatid="378" lane="2" points="432" resultid="2813" swimtime="00:00:32.31"><SPLITS/></RESULT><RESULT eventid="39" heatid="447" lane="1" points="495" resultid="3336" swimtime="00:01:05.33"><SPLITS><SPLIT distance="50" swimtime="00:00:32.17"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="603" birthdate="2015-01-01" firstname="Theresa" gender="F" lastname="Bär" license="479601"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="31" heatid="331" lane="2" points="191" resultid="2460" swimtime="00:01:51.22"><SPLITS/></RESULT><RESULT eventid="39" heatid="428" lane="2" points="186" resultid="3187" swimtime="00:01:30.51"><SPLITS><SPLIT distance="50" swimtime="00:00:43.14"/></SPLITS></RESULT></RESULTS></ATHLETE></ATHLETES><RELAYS/></CLUB><CLUB code="4562" name="TV Parsberg" nation="GER" region="02" shortname="Parsberg" type="CLUB"><CONTACT city="Lupburg" email="inesschmid.privat@t-online.de" fax="09492/902042" name="Schmid, Ines" phone="09492/902040" street="Ritter-Christoph-Weg 16" zip="92331"/><OFFICIALS/><ATHLETES><ATHLETE athleteid="23" birthdate="2013-01-01" firstname="Rosalie" gender="F" lastname="Eichenseher" license="490876"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="4" lane="3" points="115" resultid="23" swimtime="00:01:00.20"><SPLITS/></RESULT><RESULT eventid="9" heatid="105" lane="5" points="153" resultid="789" swimtime="00:00:44.25"><SPLITS/></RESULT><RESULT eventid="27" heatid="259" lane="6" points="181" resultid="1921" swimtime="00:00:47.62"><SPLITS/></RESULT><RESULT eventid="31" heatid="327" lane="2" points="134" resultid="2429" swimtime="00:02:05.26"><SPLITS><SPLIT distance="50" swimtime="00:00:57.47"/></SPLITS></RESULT><RESULT eventid="35" heatid="363" lane="1" points="67" resultid="2696" swimtime="00:01:00.13"><SPLITS/></RESULT><RESULT eventid="39" heatid="420" lane="6" points="105" resultid="3130" swimtime="00:01:49.54"><SPLITS><SPLIT distance="50" swimtime="00:00:51.47"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="128" birthdate="2012-01-01" firstname="Lena" gender="F" lastname="Pappler" license="453904"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="17" lane="4" points="310" resultid="128" swimtime="00:00:43.26"><SPLITS/></RESULT><RESULT eventid="7" heatid="89" lane="1" points="321" resultid="665" swimtime="00:03:22.75"><SPLITS><SPLIT distance="50" swimtime="00:00:45.30"/><SPLIT distance="100" swimtime="00:01:36.84"/><SPLIT distance="150" swimtime="00:02:31.99"/></SPLITS></RESULT><RESULT eventid="9" heatid="116" lane="4" points="314" resultid="876" swimtime="00:00:34.80"><SPLITS/></RESULT><RESULT eventid="27" heatid="262" lane="5" points="267" resultid="1944" swimtime="00:00:41.87"><SPLITS/></RESULT><RESULT eventid="31" heatid="338" lane="4" points="323" resultid="2518" swimtime="00:01:33.39"><SPLITS><SPLIT distance="50" swimtime="00:00:43.53"/></SPLITS></RESULT><RESULT eventid="35" heatid="369" lane="2" points="201" resultid="2744" swimtime="00:00:41.68"><SPLITS/></RESULT><RESULT eventid="39" heatid="431" lane="5" points="282" resultid="3214" swimtime="00:01:18.79"><SPLITS><SPLIT distance="50" swimtime="00:00:37.50"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="149" birthdate="2010-01-01" firstname="Anna-Lena" gender="F" lastname="Weber" license="425608"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="20" lane="1" points="358" resultid="149" swimtime="00:00:41.25"><SPLITS/></RESULT><RESULT eventid="5" heatid="66" lane="8" points="286" resultid="496" swimtime="00:01:24.12"><SPLITS><SPLIT distance="50" swimtime="00:00:38.70"/></SPLITS></RESULT><RESULT eventid="9" heatid="123" lane="7" points="385" resultid="934" swimtime="00:00:32.53"><SPLITS/></RESULT><RESULT eventid="13" heatid="204" lane="6" resultid="1549" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="27" heatid="266" lane="5" points="369" resultid="1976" swimtime="00:00:37.61"><SPLITS/></RESULT><RESULT eventid="39" heatid="444" lane="8" points="393" resultid="3320" swimtime="00:01:10.56"><SPLITS><SPLIT distance="50" swimtime="00:00:33.82"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="288" birthdate="2010-01-01" firstname="Jonas" gender="M" lastname="Pappler" license="446807"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="38" lane="6" points="377" resultid="288" swimtime="00:00:35.90"><SPLITS/></RESULT><RESULT eventid="6" heatid="74" lane="1" points="249" resultid="551" swimtime="00:01:18.57"><SPLITS><SPLIT distance="50" swimtime="00:00:32.03"/></SPLITS></RESULT><RESULT eventid="10" heatid="151" lane="6" points="439" resultid="1143" swimtime="00:00:27.50"><SPLITS/></RESULT><RESULT eventid="28" heatid="285" lane="1" points="304" resultid="2116" swimtime="00:00:35.25"><SPLITS/></RESULT><RESULT eventid="32" heatid="353" lane="5" points="323" resultid="2631" swimtime="00:01:22.84"><SPLITS><SPLIT distance="50" swimtime="00:00:36.71"/></SPLITS></RESULT><RESULT eventid="36" heatid="395" lane="2" points="356" resultid="2943" swimtime="00:00:31.42"><SPLITS/></RESULT><RESULT eventid="40" heatid="469" lane="4" resultid="3509" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="585" birthdate="2010-01-01" firstname="Anna" gender="F" lastname="Eckert" license="412523"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="27" heatid="265" lane="1" points="335" resultid="1964" swimtime="00:00:38.84"><SPLITS/></RESULT><RESULT eventid="35" heatid="368" lane="5" points="257" resultid="2739" swimtime="00:00:38.38"><SPLITS/></RESULT><RESULT eventid="39" heatid="433" lane="1" points="272" resultid="3226" swimtime="00:01:19.76"><SPLITS><SPLIT distance="50" swimtime="00:00:38.16"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="591" birthdate="2013-01-01" firstname="Thomas" gender="M" lastname="Volz" license="463742"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="28" heatid="275" lane="5" resultid="2043" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="30" heatid="310" lane="6" resultid="2309" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="32" heatid="347" lane="4" resultid="2585" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="36" heatid="383" lane="6" resultid="2855" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="40" heatid="454" lane="7" resultid="3396" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="604" birthdate="2001-01-01" firstname="Simona" gender="F" lastname="Stöckl" license="264312"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="31" heatid="342" lane="1" points="409" resultid="2547" swimtime="00:01:26.37"><SPLITS><SPLIT distance="50" swimtime="00:00:40.48"/></SPLITS></RESULT><RESULT eventid="35" heatid="380" lane="3" points="399" resultid="2830" swimtime="00:00:33.18"><SPLITS/></RESULT></RESULTS></ATHLETE></ATHLETES><RELAYS/></CLUB><CLUB code="4492" name="TSV Vaterstetten" nation="GER" region="02" shortname="Vaterstn" type="CLUB"><CONTACT city="Vaterstetten" country="GER" email="schwimmen@tsv-vaterstetten.de" name="Ostermaier, Sabine" phone="08106-6464" street="Philipp-Maas-Weg 14" zip="85591"/><OFFICIALS/><ATHLETES><ATHLETE athleteid="28" birthdate="2017-01-01" firstname="Sandra" gender="F" lastname="Hocke" license="498053"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="4" lane="8" points="86" resultid="28" swimtime="00:01:06.34"><SPLITS/></RESULT><RESULT eventid="9" heatid="105" lane="2" points="107" resultid="786" swimtime="00:00:49.79"><SPLITS/></RESULT><RESULT eventid="13" heatid="192" lane="2" points="98" resultid="1449" swimtime="00:02:04.54"><SPLITS><SPLIT distance="50" swimtime="00:01:00.34"/></SPLITS></RESULT><RESULT eventid="27" heatid="255" lane="5" points="95" resultid="1888" swimtime="00:00:59.10"><SPLITS/></RESULT><RESULT eventid="39" heatid="422" lane="3" points="80" resultid="3141" swimtime="00:01:59.82"><SPLITS><SPLIT distance="50" swimtime="00:00:53.65"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="31" birthdate="2016-01-01" firstname="Vanessa" gender="F" lastname="Wiegartner" license="482092"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="5" lane="3" points="169" resultid="31" swimtime="00:00:52.97"><SPLITS/></RESULT><RESULT eventid="9" heatid="106" lane="6" points="165" resultid="798" swimtime="00:00:43.13"><SPLITS/></RESULT><RESULT eventid="13" heatid="194" lane="3" points="169" resultid="1466" swimtime="00:01:43.87"><SPLITS><SPLIT distance="50" swimtime="00:00:49.32"/></SPLITS></RESULT><RESULT eventid="29" heatid="290" lane="7" points="152" resultid="2157" swimtime="00:03:31.39"><SPLITS><SPLIT distance="50" swimtime="00:00:47.27"/><SPLIT distance="100" swimtime="00:01:42.25"/><SPLIT distance="150" swimtime="00:02:37.71"/></SPLITS></RESULT><RESULT eventid="31" heatid="331" lane="7" points="176" resultid="2465" swimtime="00:01:54.27"><SPLITS/></RESULT><RESULT eventid="35" heatid="364" lane="6" points="83" resultid="2708" swimtime="00:00:55.92"><SPLITS/></RESULT><RESULT eventid="39" heatid="426" lane="1" points="128" resultid="3170" swimtime="00:01:42.38"><SPLITS><SPLIT distance="50" swimtime="00:00:48.95"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="41" birthdate="2015-01-01" firstname="Franziska" gender="F" lastname="Krenz" license="488394"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="6" lane="5" points="172" resultid="41" swimtime="00:00:52.68"><SPLITS/></RESULT><RESULT eventid="9" heatid="104" lane="5" points="157" resultid="781" swimtime="00:00:43.84"><SPLITS/></RESULT><RESULT eventid="13" heatid="194" lane="6" points="156" resultid="1469" swimtime="00:01:46.54"><SPLITS><SPLIT distance="50" swimtime="00:00:51.63"/></SPLITS></RESULT><RESULT eventid="27" heatid="257" lane="5" points="159" resultid="1904" swimtime="00:00:49.74"><SPLITS/></RESULT><RESULT eventid="29" heatid="289" lane="8" points="143" resultid="2150" swimtime="00:03:35.89"><SPLITS><SPLIT distance="50" swimtime="00:00:49.68"/><SPLIT distance="100" swimtime="00:01:44.90"/><SPLIT distance="150" swimtime="00:02:44.21"/></SPLITS></RESULT><RESULT eventid="37" heatid="402" lane="7" points="165" resultid="2998" swimtime="00:03:44.63"><SPLITS><SPLIT distance="50" swimtime="00:00:54.11"/><SPLIT distance="100" swimtime="00:01:51.95"/><SPLIT distance="150" swimtime="00:02:50.12"/></SPLITS></RESULT><RESULT eventid="39" heatid="427" lane="8" points="139" resultid="3185" swimtime="00:01:39.68"><SPLITS><SPLIT distance="50" swimtime="00:00:47.65"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="43" birthdate="2016-01-01" firstname="Ella" gender="F" lastname="Oettrich" license="482090"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="6" lane="7" points="142" resultid="43" swimtime="00:00:56.14"><SPLITS/></RESULT><RESULT eventid="9" heatid="106" lane="7" points="193" resultid="799" swimtime="00:00:40.91"><SPLITS/></RESULT><RESULT eventid="13" heatid="196" lane="1" points="187" resultid="1480" swimtime="00:01:40.41"><SPLITS><SPLIT distance="50" swimtime="00:00:47.86"/></SPLITS></RESULT><RESULT eventid="27" heatid="259" lane="8" points="212" resultid="1923" swimtime="00:00:45.23"><SPLITS/></RESULT><RESULT eventid="29" heatid="290" lane="2" points="150" resultid="2152" swimtime="00:03:32.62"><SPLITS><SPLIT distance="50" swimtime="00:00:47.77"/><SPLIT distance="100" swimtime="00:01:44.33"/><SPLIT distance="150" swimtime="00:02:39.91"/></SPLITS></RESULT><RESULT eventid="37" heatid="402" lane="6" points="191" resultid="2997" swimtime="00:03:34.08"><SPLITS><SPLIT distance="100" swimtime="00:01:46.16"/></SPLITS></RESULT><RESULT eventid="39" heatid="426" lane="7" points="140" resultid="3176" swimtime="00:01:39.57"><SPLITS><SPLIT distance="50" swimtime="00:00:45.13"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="48" birthdate="2015-01-01" firstname="Xinchen" gender="F" lastname="Du" license="482658"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="7" lane="4" points="151" resultid="48" swimtime="00:00:55.00"><SPLITS/></RESULT><RESULT eventid="9" heatid="109" lane="1" points="150" resultid="817" swimtime="00:00:44.46"><SPLITS/></RESULT><RESULT eventid="13" heatid="194" lane="7" points="136" resultid="1470" swimtime="00:01:51.71"><SPLITS><SPLIT distance="50" swimtime="00:00:53.63"/></SPLITS></RESULT><RESULT eventid="27" heatid="258" lane="8" points="135" resultid="1915" swimtime="00:00:52.47"><SPLITS/></RESULT><RESULT eventid="31" heatid="330" lane="8" points="148" resultid="2458" swimtime="00:02:01.12"><SPLITS/></RESULT><RESULT eventid="39" heatid="423" lane="3" points="141" resultid="3149" swimtime="00:01:39.30"><SPLITS><SPLIT distance="50" swimtime="00:00:46.09"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="54" birthdate="2014-01-01" firstname="Emily" gender="F" lastname="O'Connell" license="460786"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="8" lane="2" points="169" resultid="54" swimtime="00:00:52.91"><SPLITS/></RESULT><RESULT eventid="11" heatid="160" lane="2" points="194" resultid="1204" swimtime="00:03:37.86"><SPLITS><SPLIT distance="50" swimtime="00:00:51.80"/><SPLIT distance="100" swimtime="00:01:40.88"/><SPLIT distance="150" swimtime="00:02:42.55"/></SPLITS></RESULT><RESULT eventid="13" heatid="198" lane="4" points="245" resultid="1499" swimtime="00:01:31.77"><SPLITS><SPLIT distance="50" swimtime="00:00:44.52"/></SPLITS></RESULT><RESULT eventid="27" heatid="261" lane="6" points="270" resultid="1937" swimtime="00:00:41.74"><SPLITS/></RESULT><RESULT eventid="29" heatid="289" lane="5" points="171" resultid="2147" swimtime="00:03:23.41"><SPLITS><SPLIT distance="50" swimtime="00:00:46.21"/><SPLIT distance="100" swimtime="00:01:39.23"/><SPLIT distance="150" swimtime="00:02:32.24"/></SPLITS></RESULT><RESULT eventid="37" heatid="403" lane="4" points="237" resultid="3002" swimtime="00:03:19.19"><SPLITS><SPLIT distance="50" swimtime="00:00:46.16"/><SPLIT distance="100" swimtime="00:01:37.45"/><SPLIT distance="150" swimtime="00:02:30.02"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="56" birthdate="2014-01-01" firstname="Charlotte" gender="F" lastname="Gerhardt" license="460781"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="8" lane="4" points="209" resultid="56" swimtime="00:00:49.37"><SPLITS/></RESULT><RESULT eventid="7" heatid="83" lane="3" points="219" resultid="620" swimtime="00:03:50.21"><SPLITS><SPLIT distance="50" swimtime="00:00:51.82"/><SPLIT distance="100" swimtime="00:01:52.99"/><SPLIT distance="150" swimtime="00:02:52.31"/></SPLITS></RESULT><RESULT eventid="9" heatid="112" lane="3" points="273" resultid="843" swimtime="00:00:36.45"><SPLITS/></RESULT><RESULT eventid="11" heatid="161" lane="6" points="257" resultid="1216" swimtime="00:03:18.22"><SPLITS><SPLIT distance="50" swimtime="00:00:45.17"/><SPLIT distance="100" swimtime="00:01:36.61"/><SPLIT distance="150" swimtime="00:02:36.07"/></SPLITS></RESULT><RESULT eventid="29" heatid="294" lane="5" points="259" resultid="2186" swimtime="00:02:57.08"><SPLITS><SPLIT distance="50" swimtime="00:00:39.30"/><SPLIT distance="100" swimtime="00:01:25.57"/><SPLIT distance="150" swimtime="00:02:13.56"/></SPLITS></RESULT><RESULT eventid="31" heatid="334" lane="4" points="207" resultid="2486" swimtime="00:01:48.25"><SPLITS><SPLIT distance="50" swimtime="00:00:50.10"/></SPLITS></RESULT><RESULT eventid="39" heatid="431" lane="6" points="267" resultid="3215" swimtime="00:01:20.23"><SPLITS><SPLIT distance="50" swimtime="00:00:37.18"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="69" birthdate="2015-01-01" firstname="Carla" gender="F" lastname="May" license="465838"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="10" lane="1" points="175" resultid="69" swimtime="00:00:52.38"><SPLITS/></RESULT><RESULT eventid="7" heatid="82" lane="8" points="177" resultid="617" swimtime="00:04:07.13"><SPLITS><SPLIT distance="50" swimtime="00:00:56.98"/><SPLIT distance="100" swimtime="00:01:58.47"/><SPLIT distance="150" swimtime="00:03:05.12"/></SPLITS></RESULT><RESULT eventid="9" heatid="106" lane="1" points="163" resultid="793" swimtime="00:00:43.32"><SPLITS/></RESULT><RESULT eventid="13" heatid="193" lane="5" points="155" resultid="1460" swimtime="00:01:46.79"><SPLITS/></RESULT><RESULT eventid="29" heatid="288" lane="3" points="137" resultid="2139" swimtime="00:03:38.63"><SPLITS><SPLIT distance="50" swimtime="00:00:49.30"/><SPLIT distance="100" swimtime="00:01:43.82"/><SPLIT distance="150" swimtime="00:02:43.34"/></SPLITS></RESULT><RESULT eventid="31" heatid="331" lane="4" points="172" resultid="2462" swimtime="00:01:55.30"><SPLITS/></RESULT><RESULT eventid="39" heatid="423" lane="5" points="140" resultid="3151" swimtime="00:01:39.37"><SPLITS><SPLIT distance="50" swimtime="00:00:46.46"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="74" birthdate="2015-01-01" firstname="Julia" gender="F" lastname="Hocke" license="464715"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="10" lane="6" points="174" resultid="74" swimtime="00:00:52.47"><SPLITS/></RESULT><RESULT eventid="7" heatid="82" lane="1" points="180" resultid="610" swimtime="00:04:05.85"><SPLITS><SPLIT distance="50" swimtime="00:00:56.49"/><SPLIT distance="100" swimtime="00:01:59.90"/><SPLIT distance="150" swimtime="00:03:05.39"/></SPLITS></RESULT><RESULT eventid="9" heatid="108" lane="7" points="168" resultid="815" swimtime="00:00:42.86"><SPLITS/></RESULT><RESULT eventid="13" heatid="195" lane="8" points="151" resultid="1479" swimtime="00:01:47.66"><SPLITS><SPLIT distance="50" swimtime="00:00:52.44"/></SPLITS></RESULT><RESULT eventid="27" heatid="259" lane="3" points="155" resultid="1918" swimtime="00:00:50.21"><SPLITS/></RESULT><RESULT eventid="29" heatid="288" lane="4" points="123" resultid="2140" swimtime="00:03:46.61"><SPLITS><SPLIT distance="50" swimtime="00:00:49.25"/><SPLIT distance="100" swimtime="00:01:49.21"/><SPLIT distance="150" swimtime="00:02:47.99"/></SPLITS></RESULT><RESULT eventid="37" heatid="402" lane="1" points="152" resultid="2992" swimtime="00:03:50.97"><SPLITS><SPLIT distance="50" swimtime="00:00:54.55"/><SPLIT distance="100" swimtime="00:01:53.84"/><SPLIT distance="150" swimtime="00:02:56.10"/></SPLITS></RESULT><RESULT eventid="39" heatid="426" lane="2" points="125" resultid="3171" swimtime="00:01:43.33"><SPLITS><SPLIT distance="50" swimtime="00:00:48.13"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="82" birthdate="2014-01-01" firstname="Orla" gender="F" lastname="O'Connell" license="460787"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="11" lane="6" points="193" resultid="82" swimtime="00:00:50.63"><SPLITS/></RESULT><RESULT eventid="7" heatid="82" lane="7" points="198" resultid="616" swimtime="00:03:58.29"><SPLITS><SPLIT distance="50" swimtime="00:00:54.21"/><SPLIT distance="100" swimtime="00:01:55.19"/><SPLIT distance="150" swimtime="00:02:57.04"/></SPLITS></RESULT><RESULT eventid="13" heatid="195" lane="1" points="187" resultid="1472" swimtime="00:01:40.29"><SPLITS><SPLIT distance="50" swimtime="00:00:47.03"/></SPLITS></RESULT><RESULT eventid="29" heatid="289" lane="2" points="155" resultid="2144" swimtime="00:03:30.08"><SPLITS><SPLIT distance="50" swimtime="00:00:45.88"/><SPLIT distance="100" swimtime="00:01:40.27"/><SPLIT distance="150" swimtime="00:02:36.01"/></SPLITS></RESULT><RESULT eventid="31" heatid="333" lane="2" points="196" resultid="2476" swimtime="00:01:50.37"><SPLITS><SPLIT distance="50" swimtime="00:00:52.67"/></SPLITS></RESULT><RESULT eventid="39" heatid="425" lane="7" points="165" resultid="3168" swimtime="00:01:34.20"><SPLITS><SPLIT distance="50" swimtime="00:00:43.86"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="89" birthdate="2014-01-01" firstname="Antonia" gender="F" lastname="Resch" license="465839"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="12" lane="5" points="188" resultid="89" swimtime="00:00:51.14"><SPLITS/></RESULT><RESULT eventid="7" heatid="82" lane="2" points="229" resultid="611" swimtime="00:03:46.93"><SPLITS><SPLIT distance="50" swimtime="00:00:54.07"/><SPLIT distance="100" swimtime="00:01:52.58"/><SPLIT distance="150" swimtime="00:02:50.72"/></SPLITS></RESULT><RESULT eventid="9" heatid="110" lane="7" points="190" resultid="831" swimtime="00:00:41.12"><SPLITS/></RESULT><RESULT eventid="29" heatid="290" lane="1" points="164" resultid="2151" swimtime="00:03:26.25"><SPLITS><SPLIT distance="50" swimtime="00:00:44.32"/><SPLIT distance="100" swimtime="00:01:37.32"/><SPLIT distance="150" swimtime="00:02:32.49"/></SPLITS></RESULT><RESULT eventid="31" heatid="334" lane="7" points="191" resultid="2489" swimtime="00:01:51.27"><SPLITS><SPLIT distance="50" swimtime="00:00:53.17"/></SPLITS></RESULT><RESULT eventid="39" heatid="425" lane="8" points="168" resultid="3169" swimtime="00:01:33.64"><SPLITS><SPLIT distance="50" swimtime="00:00:45.99"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="96" birthdate="2014-01-01" firstname="Jule" gender="F" lastname="Ostermaier" license="455479"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="13" lane="4" points="236" resultid="96" swimtime="00:00:47.39"><SPLITS/></RESULT><RESULT eventid="7" heatid="82" lane="6" points="258" resultid="615" swimtime="00:03:38.07"><SPLITS><SPLIT distance="50" swimtime="00:00:50.24"/><SPLIT distance="100" swimtime="00:01:46.11"/><SPLIT distance="150" swimtime="00:02:42.68"/></SPLITS></RESULT><RESULT eventid="11" heatid="160" lane="3" points="258" resultid="1205" swimtime="00:03:17.91"><SPLITS><SPLIT distance="50" swimtime="00:00:45.46"/><SPLIT distance="100" swimtime="00:01:34.98"/><SPLIT distance="150" swimtime="00:02:32.11"/></SPLITS></RESULT><RESULT eventid="29" heatid="292" lane="4" points="265" resultid="2169" swimtime="00:02:55.82"><SPLITS><SPLIT distance="50" swimtime="00:00:39.37"/><SPLIT distance="100" swimtime="00:01:24.01"/><SPLIT distance="150" swimtime="00:02:10.46"/></SPLITS></RESULT><RESULT eventid="37" heatid="403" lane="8" points="238" resultid="3006" swimtime="00:03:18.83"><SPLITS><SPLIT distance="50" swimtime="00:00:47.75"/><SPLIT distance="100" swimtime="00:01:37.10"/><SPLIT distance="150" swimtime="00:02:30.50"/></SPLITS></RESULT><RESULT eventid="39" heatid="431" lane="1" points="235" resultid="3210" swimtime="00:01:23.72"><SPLITS><SPLIT distance="50" swimtime="00:00:39.42"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="97" birthdate="2015-01-01" firstname="Greta" gender="F" lastname="Kaltenbrunner" license="465024"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="13" lane="5" points="220" resultid="97" swimtime="00:00:48.49"><SPLITS/></RESULT><RESULT eventid="7" heatid="83" lane="4" points="211" resultid="621" swimtime="00:03:53.13"><SPLITS><SPLIT distance="50" swimtime="00:00:51.59"/><SPLIT distance="100" swimtime="00:01:52.24"/><SPLIT distance="150" swimtime="00:02:53.48"/></SPLITS></RESULT><RESULT eventid="9" heatid="109" lane="8" points="145" resultid="824" swimtime="00:00:44.96"><SPLITS/></RESULT><RESULT eventid="13" heatid="193" lane="8" points="150" resultid="1463" swimtime="00:01:48.05"><SPLITS><SPLIT distance="50" swimtime="00:00:52.58"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="107" birthdate="2014-01-01" firstname="Johanna" gender="F" lastname="Rinderknecht" license="443249"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="14" lane="7" points="243" resultid="107" swimtime="00:00:46.89"><SPLITS/></RESULT><RESULT eventid="7" heatid="83" lane="5" points="229" resultid="622" swimtime="00:03:46.98"><SPLITS><SPLIT distance="50" swimtime="00:00:52.61"/><SPLIT distance="100" swimtime="00:01:51.72"/><SPLIT distance="150" swimtime="00:02:50.60"/></SPLITS></RESULT><RESULT eventid="9" heatid="110" lane="8" points="230" resultid="832" swimtime="00:00:38.59"><SPLITS/></RESULT><RESULT eventid="29" heatid="293" lane="1" points="217" resultid="2174" swimtime="00:03:07.90"><SPLITS><SPLIT distance="50" swimtime="00:00:43.05"/><SPLIT distance="100" swimtime="00:01:30.36"/><SPLIT distance="150" swimtime="00:02:21.40"/></SPLITS></RESULT><RESULT eventid="31" heatid="334" lane="5" points="241" resultid="2487" swimtime="00:01:43.02"><SPLITS><SPLIT distance="50" swimtime="00:00:48.37"/></SPLITS></RESULT><RESULT eventid="39" heatid="429" lane="6" points="234" resultid="3199" swimtime="00:01:23.84"><SPLITS><SPLIT distance="50" swimtime="00:00:39.42"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="169" birthdate="2009-01-01" firstname="Isabelle" gender="F" lastname="O'Connell" license="415011"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="22" lane="7" points="464" resultid="169" swimtime="00:00:37.84"><SPLITS/></RESULT><RESULT eventid="7" heatid="90" lane="1" points="447" resultid="673" swimtime="00:03:01.69"><SPLITS><SPLIT distance="50" swimtime="00:00:42.39"/><SPLIT distance="100" swimtime="00:01:28.32"/><SPLIT distance="150" swimtime="00:02:17.31"/></SPLITS></RESULT><RESULT eventid="9" heatid="121" lane="7" points="450" resultid="918" swimtime="00:00:30.87"><SPLITS/></RESULT><RESULT eventid="11" heatid="170" lane="1" points="411" resultid="1283" swimtime="00:02:49.60"><SPLITS><SPLIT distance="50" swimtime="00:00:38.23"/><SPLIT distance="100" swimtime="00:01:19.50"/><SPLIT distance="150" swimtime="00:02:10.10"/></SPLITS></RESULT><RESULT eventid="27" heatid="265" lane="3" points="397" resultid="1966" swimtime="00:00:36.68"><SPLITS/></RESULT><RESULT eventid="31" heatid="342" lane="6" points="463" resultid="2552" swimtime="00:01:22.84"><SPLITS><SPLIT distance="50" swimtime="00:00:39.38"/></SPLITS></RESULT><RESULT eventid="39" heatid="440" lane="5" points="431" resultid="3285" swimtime="00:01:08.43"><SPLITS><SPLIT distance="50" swimtime="00:00:32.57"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="177" birthdate="2012-01-01" firstname="Lena" gender="F" lastname="Ostermaier" license="436077"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="23" lane="7" points="501" resultid="177" swimtime="00:00:36.89"><SPLITS/></RESULT><RESULT eventid="5" heatid="69" lane="1" points="329" resultid="512" swimtime="00:01:20.35"><SPLITS><SPLIT distance="50" swimtime="00:00:37.25"/></SPLITS></RESULT><RESULT eventid="11" heatid="171" lane="3" points="468" resultid="1293" swimtime="00:02:42.43"><SPLITS><SPLIT distance="50" swimtime="00:00:35.08"/><SPLIT distance="100" swimtime="00:01:17.28"/><SPLIT distance="150" swimtime="00:02:05.17"/></SPLITS></RESULT><RESULT eventid="27" heatid="266" lane="2" points="380" resultid="1973" swimtime="00:00:37.22"><SPLITS/></RESULT><RESULT eventid="31" heatid="343" lane="2" points="499" resultid="2556" swimtime="00:01:20.84"><SPLITS><SPLIT distance="50" swimtime="00:00:39.36"/></SPLITS></RESULT><RESULT eventid="35" heatid="378" lane="7" points="381" resultid="2818" swimtime="00:00:33.69"><SPLITS/></RESULT><RESULT eventid="39" heatid="441" lane="4" points="435" resultid="3292" swimtime="00:01:08.21"><SPLITS><SPLIT distance="50" swimtime="00:00:32.27"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="178" birthdate="2004-01-01" firstname="Marlen Seraphine" gender="F" lastname="Görlach" license="306532"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="23" lane="8" points="393" resultid="178" swimtime="00:00:40.00"><SPLITS/></RESULT><RESULT eventid="5" heatid="70" lane="2" points="426" resultid="521" swimtime="00:01:13.73"><SPLITS><SPLIT distance="50" swimtime="00:00:33.94"/></SPLITS></RESULT><RESULT eventid="9" heatid="130" lane="8" points="441" resultid="989" swimtime="00:00:31.08"><SPLITS/></RESULT><RESULT eventid="11" heatid="173" lane="6" points="446" resultid="1312" swimtime="00:02:44.99"><SPLITS><SPLIT distance="50" swimtime="00:00:34.64"/><SPLIT distance="100" swimtime="00:01:18.19"/><SPLIT distance="150" swimtime="00:02:06.25"/></SPLITS></RESULT><RESULT eventid="29" heatid="306" lane="6" points="461" resultid="2280" swimtime="00:02:26.17"><SPLITS><SPLIT distance="50" swimtime="00:00:32.92"/><SPLIT distance="100" swimtime="00:01:09.49"/><SPLIT distance="150" swimtime="00:01:47.04"/></SPLITS></RESULT><RESULT eventid="35" heatid="381" lane="3" points="431" resultid="2838" swimtime="00:00:32.32"><SPLITS/></RESULT><RESULT eventid="39" heatid="449" lane="3" points="521" resultid="3353" swimtime="00:01:04.23"><SPLITS><SPLIT distance="50" swimtime="00:00:31.04"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="206" birthdate="2015-01-01" firstname="Finn" gender="M" lastname="Arnold" license="465023"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="28" lane="2" points="105" resultid="206" swimtime="00:00:54.95"><SPLITS/></RESULT><RESULT eventid="10" heatid="138" lane="7" points="134" resultid="1042" swimtime="00:00:40.79"><SPLITS/></RESULT><RESULT eventid="14" heatid="214" lane="7" points="104" resultid="1627" swimtime="00:01:49.65"><SPLITS><SPLIT distance="50" swimtime="00:00:51.62"/></SPLITS></RESULT><RESULT eventid="28" heatid="278" lane="1" points="99" resultid="2061" swimtime="00:00:51.16"><SPLITS/></RESULT><RESULT eventid="30" heatid="311" lane="7" points="107" resultid="2317" swimtime="00:03:34.56"><SPLITS><SPLIT distance="50" swimtime="00:00:48.30"/><SPLIT distance="100" swimtime="00:01:46.00"/><SPLIT distance="150" swimtime="00:02:42.11"/></SPLITS></RESULT><RESULT eventid="38" heatid="414" lane="1" points="88" resultid="3083" swimtime="00:04:11.45"><SPLITS><SPLIT distance="50" swimtime="00:00:57.46"/><SPLIT distance="100" swimtime="00:02:03.23"/><SPLIT distance="150" swimtime="00:03:08.74"/></SPLITS></RESULT><RESULT eventid="40" heatid="456" lane="7" resultid="3411" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="220" birthdate="2014-01-01" firstname="Jan" gender="M" lastname="Rathmann" license="460792"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="29" lane="8" points="102" resultid="220" swimtime="00:00:55.46"><SPLITS/></RESULT><RESULT eventid="10" heatid="137" lane="6" points="155" resultid="1034" swimtime="00:00:38.89"><SPLITS/></RESULT><RESULT eventid="14" heatid="212" lane="6" points="104" resultid="1610" swimtime="00:01:49.45"><SPLITS><SPLIT distance="50" swimtime="00:00:52.45"/></SPLITS></RESULT><RESULT eventid="28" heatid="276" lane="5" points="115" resultid="2051" swimtime="00:00:48.65"><SPLITS/></RESULT><RESULT eventid="30" heatid="310" lane="2" points="110" resultid="2305" swimtime="00:03:32.64"><SPLITS><SPLIT distance="50" swimtime="00:00:47.51"/><SPLIT distance="100" swimtime="00:01:42.62"/><SPLIT distance="150" swimtime="00:02:39.91"/></SPLITS></RESULT><RESULT eventid="40" heatid="454" lane="1" points="130" resultid="3390" swimtime="00:01:32.37"><SPLITS><SPLIT distance="50" swimtime="00:00:43.35"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="236" birthdate="2015-01-01" firstname="Fjonn" gender="M" lastname="Bartel" license="488385"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="31" lane="8" points="131" resultid="236" swimtime="00:00:51.05"><SPLITS/></RESULT><RESULT eventid="8" heatid="93" lane="6" points="149" resultid="702" swimtime="00:03:57.29"><SPLITS><SPLIT distance="50" swimtime="00:00:53.32"/><SPLIT distance="100" swimtime="00:01:54.02"/><SPLIT distance="150" swimtime="00:02:56.12"/></SPLITS></RESULT><RESULT eventid="10" heatid="135" lane="1" points="113" resultid="1013" swimtime="00:00:43.16"><SPLITS/></RESULT><RESULT eventid="14" heatid="213" lane="4" points="123" resultid="1616" swimtime="00:01:43.62"><SPLITS><SPLIT distance="50" swimtime="00:00:49.07"/></SPLITS></RESULT><RESULT eventid="30" heatid="311" lane="8" points="124" resultid="2318" swimtime="00:03:24.31"><SPLITS><SPLIT distance="50" swimtime="00:00:47.59"/><SPLIT distance="100" swimtime="00:01:39.43"/><SPLIT distance="150" swimtime="00:02:33.88"/></SPLITS></RESULT><RESULT eventid="32" heatid="347" lane="1" points="116" resultid="2582" swimtime="00:01:56.50"><SPLITS><SPLIT distance="50" swimtime="00:00:56.46"/></SPLITS></RESULT><RESULT eventid="40" heatid="454" lane="4" points="117" resultid="3393" swimtime="00:01:35.60"><SPLITS><SPLIT distance="50" swimtime="00:00:45.74"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="261" birthdate="2012-01-01" firstname="Vitus" gender="M" lastname="Werler" license="441354"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="35" lane="3" points="216" resultid="261" swimtime="00:00:43.21"><SPLITS/></RESULT><RESULT eventid="8" heatid="97" lane="4" points="240" resultid="729" swimtime="00:03:22.46"><SPLITS><SPLIT distance="50" swimtime="00:00:42.79"/><SPLIT distance="100" swimtime="00:01:36.23"/><SPLIT distance="150" swimtime="00:02:30.67"/></SPLITS></RESULT><RESULT comment="16:21 Der Sportler hat die Teilstrecke Rücken nicht in Rückenlage beendet" eventid="12" heatid="180" lane="7" resultid="1364" status="DSQ" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="32" heatid="351" lane="3" points="254" resultid="2614" swimtime="00:01:29.80"><SPLITS><SPLIT distance="50" swimtime="00:00:42.29"/></SPLITS></RESULT><RESULT eventid="36" heatid="390" lane="7" points="171" resultid="2908" swimtime="00:00:40.08"><SPLITS/></RESULT><RESULT eventid="40" heatid="463" lane="1" points="267" resultid="3460" swimtime="00:01:12.70"><SPLITS><SPLIT distance="50" swimtime="00:00:35.38"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="275" birthdate="2010-01-01" firstname="Luca" gender="M" lastname="Liguori" license="415014"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="37" lane="1" points="380" resultid="275" swimtime="00:00:35.80"><SPLITS/></RESULT><RESULT eventid="8" heatid="99" lane="7" points="348" resultid="747" swimtime="00:02:58.94"><SPLITS><SPLIT distance="50" swimtime="00:00:39.84"/><SPLIT distance="100" swimtime="00:01:27.40"/><SPLIT distance="150" swimtime="00:02:14.24"/></SPLITS></RESULT><RESULT eventid="10" heatid="147" lane="4" points="400" resultid="1109" swimtime="00:00:28.37"><SPLITS/></RESULT><RESULT eventid="14" heatid="221" lane="1" points="262" resultid="1674" swimtime="00:01:20.56"><SPLITS><SPLIT distance="50" swimtime="00:00:40.74"/></SPLITS></RESULT><RESULT eventid="28" heatid="283" lane="5" points="296" resultid="2105" swimtime="00:00:35.57"><SPLITS/></RESULT><RESULT eventid="32" heatid="353" lane="7" points="403" resultid="2633" swimtime="00:01:16.95"><SPLITS><SPLIT distance="50" swimtime="00:00:35.20"/></SPLITS></RESULT><RESULT eventid="36" heatid="391" lane="7" points="275" resultid="2916" swimtime="00:00:34.24"><SPLITS/></RESULT><RESULT eventid="40" heatid="467" lane="8" points="344" resultid="3497" swimtime="00:01:06.82"><SPLITS><SPLIT distance="50" swimtime="00:00:31.07"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="296" birthdate="1998-01-01" firstname="Florian" gender="M" lastname="Maurer" license="180742"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="39" lane="6" points="469" resultid="296" swimtime="00:00:33.39"><SPLITS/></RESULT><RESULT eventid="10" heatid="152" lane="4" points="467" resultid="1149" swimtime="00:00:26.95"><SPLITS/></RESULT><RESULT eventid="12" heatid="188" lane="5" points="440" resultid="1424" swimtime="00:02:29.88"><SPLITS><SPLIT distance="50" swimtime="00:00:31.49"/><SPLIT distance="100" swimtime="00:01:12.38"/><SPLIT distance="150" swimtime="00:01:54.33"/></SPLITS></RESULT><RESULT eventid="32" heatid="355" lane="4" points="443" resultid="2645" swimtime="00:01:14.57"><SPLITS><SPLIT distance="50" swimtime="00:00:34.82"/></SPLITS></RESULT><RESULT eventid="36" heatid="397" lane="6" points="425" resultid="2963" swimtime="00:00:29.60"><SPLITS/></RESULT><RESULT eventid="40" heatid="473" lane="8" points="513" resultid="3544" swimtime="00:00:58.53"><SPLITS><SPLIT distance="50" swimtime="00:00:28.65"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="315" birthdate="2014-01-01" firstname="Paula" gender="F" lastname="Orth" license="464756"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="42" lane="6" points="242" resultid="317" swimtime="00:06:18.91"><SPLITS><SPLIT distance="100" swimtime="00:01:34.06"/><SPLIT distance="200" swimtime="00:03:09.94"/><SPLIT distance="300" swimtime="00:04:47.31"/></SPLITS></RESULT><RESULT eventid="11" heatid="162" lane="2" points="264" resultid="1220" swimtime="00:03:16.38"><SPLITS><SPLIT distance="50" swimtime="00:00:43.78"/><SPLIT distance="100" swimtime="00:01:31.71"/><SPLIT distance="150" swimtime="00:02:34.30"/></SPLITS></RESULT><RESULT eventid="13" heatid="199" lane="4" points="281" resultid="1507" swimtime="00:01:27.63"><SPLITS><SPLIT distance="50" swimtime="00:00:41.61"/></SPLITS></RESULT><RESULT eventid="19" heatid="235" lane="7" resultid="1768" swimtime="00:00:50.68"><SPLITS/></RESULT><RESULT eventid="29" heatid="294" lane="3" points="261" resultid="2184" swimtime="00:02:56.65"><SPLITS><SPLIT distance="50" swimtime="00:00:39.51"/><SPLIT distance="100" swimtime="00:01:24.84"/><SPLIT distance="150" swimtime="00:02:13.00"/></SPLITS></RESULT><RESULT eventid="37" heatid="405" lane="6" points="287" resultid="3020" swimtime="00:03:06.85"><SPLITS><SPLIT distance="50" swimtime="00:00:42.98"/><SPLIT distance="100" swimtime="00:01:31.08"/><SPLIT distance="150" swimtime="00:02:20.23"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="316" birthdate="2011-01-01" firstname="Sylvie" gender="F" lastname="Brixel" license="427026"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="42" lane="8" points="295" resultid="319" swimtime="00:05:54.93"><SPLITS><SPLIT distance="100" swimtime="00:01:24.00"/><SPLIT distance="200" swimtime="00:02:56.83"/><SPLIT distance="300" swimtime="00:04:28.47"/></SPLITS></RESULT><RESULT eventid="9" heatid="116" lane="8" points="393" resultid="880" swimtime="00:00:32.29"><SPLITS/></RESULT><RESULT eventid="13" heatid="200" lane="5" points="335" resultid="1516" swimtime="00:01:22.65"><SPLITS><SPLIT distance="50" swimtime="00:00:40.27"/></SPLITS></RESULT><RESULT eventid="27" heatid="262" lane="7" points="304" resultid="1946" swimtime="00:00:40.12"><SPLITS/></RESULT><RESULT eventid="29" heatid="298" lane="1" points="353" resultid="2214" swimtime="00:02:39.85"><SPLITS><SPLIT distance="50" swimtime="00:00:36.80"/><SPLIT distance="100" swimtime="00:01:16.91"/><SPLIT distance="150" swimtime="00:01:59.79"/></SPLITS></RESULT><RESULT eventid="35" heatid="370" lane="2" points="354" resultid="2752" swimtime="00:00:34.53"><SPLITS/></RESULT><RESULT eventid="39" heatid="438" lane="3" points="410" resultid="3268" swimtime="00:01:09.55"><SPLITS><SPLIT distance="50" swimtime="00:00:33.37"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="318" birthdate="2015-01-01" firstname="Philomena" gender="F" lastname="Werler" license="465845"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="43" lane="2" points="244" resultid="321" swimtime="00:06:17.85"><SPLITS><SPLIT distance="100" swimtime="00:01:27.60"/><SPLIT distance="200" swimtime="00:03:05.25"/><SPLIT distance="300" swimtime="00:04:42.74"/></SPLITS></RESULT><RESULT eventid="11" heatid="163" lane="6" points="264" resultid="1232" swimtime="00:03:16.53"><SPLITS><SPLIT distance="50" swimtime="00:00:44.08"/><SPLIT distance="100" swimtime="00:01:31.90"/><SPLIT distance="150" swimtime="00:02:31.66"/></SPLITS></RESULT><RESULT eventid="13" heatid="200" lane="8" points="266" resultid="1519" swimtime="00:01:29.23"><SPLITS><SPLIT distance="50" swimtime="00:00:44.49"/></SPLITS></RESULT><RESULT eventid="29" heatid="297" lane="8" points="248" resultid="2213" swimtime="00:02:59.66"><SPLITS><SPLIT distance="50" swimtime="00:00:39.82"/><SPLIT distance="100" swimtime="00:01:23.99"/><SPLIT distance="150" swimtime="00:02:13.67"/></SPLITS></RESULT><RESULT eventid="37" heatid="405" lane="1" points="274" resultid="3015" swimtime="00:03:09.69"><SPLITS><SPLIT distance="50" swimtime="00:00:45.57"/><SPLIT distance="100" swimtime="00:01:33.26"/><SPLIT distance="150" swimtime="00:02:22.87"/></SPLITS></RESULT><RESULT eventid="39" heatid="433" lane="8" points="262" resultid="3233" swimtime="00:01:20.75"><SPLITS><SPLIT distance="50" swimtime="00:00:38.89"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="319" birthdate="2013-01-01" firstname="Yara" gender="F" lastname="Gutmann" license="455400"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="43" lane="3" resultid="322" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="5" heatid="64" lane="3" resultid="475" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="9" heatid="111" lane="4" resultid="836" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="13" heatid="199" lane="6" resultid="1509" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="325" birthdate="2014-01-01" firstname="Emily" gender="F" lastname="Strasser" license="460789"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="44" lane="4" points="335" resultid="331" swimtime="00:05:40.30"><SPLITS><SPLIT distance="100" swimtime="00:01:22.17"/><SPLIT distance="200" swimtime="00:02:49.73"/><SPLIT distance="300" swimtime="00:04:17.13"/></SPLITS></RESULT><RESULT eventid="11" heatid="166" lane="2" points="331" resultid="1252" swimtime="00:03:02.30"><SPLITS><SPLIT distance="50" swimtime="00:00:40.95"/><SPLIT distance="100" swimtime="00:01:26.06"/><SPLIT distance="150" swimtime="00:02:24.02"/></SPLITS></RESULT><RESULT eventid="13" heatid="203" lane="3" points="346" resultid="1538" swimtime="00:01:21.76"><SPLITS><SPLIT distance="50" swimtime="00:00:40.02"/></SPLITS></RESULT><RESULT eventid="19" heatid="235" lane="2" resultid="1763" swimtime="00:00:51.15"><SPLITS/></RESULT><RESULT eventid="27" heatid="267" lane="1" points="329" resultid="1980" swimtime="00:00:39.07"><SPLITS/></RESULT><RESULT eventid="37" heatid="406" lane="4" points="373" resultid="3026" swimtime="00:02:51.21"><SPLITS><SPLIT distance="50" swimtime="00:00:40.15"/><SPLIT distance="100" swimtime="00:01:23.93"/><SPLIT distance="150" swimtime="00:02:08.01"/></SPLITS></RESULT><RESULT eventid="39" heatid="435" lane="3" points="351" resultid="3244" swimtime="00:01:13.30"><SPLITS><SPLIT distance="50" swimtime="00:00:35.48"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="359" birthdate="2010-01-01" firstname="Sophia" gender="F" lastname="Hofmann" license="415008"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="50" lane="4" points="440" resultid="378" swimtime="00:05:10.80"><SPLITS><SPLIT distance="100" swimtime="00:01:12.22"/><SPLIT distance="200" swimtime="00:02:32.09"/><SPLIT distance="300" swimtime="00:03:51.94"/></SPLITS></RESULT><RESULT eventid="9" heatid="125" lane="1" points="406" resultid="944" swimtime="00:00:31.94"><SPLITS/></RESULT><RESULT eventid="13" heatid="207" lane="2" points="466" resultid="1569" swimtime="00:01:14.07"><SPLITS><SPLIT distance="50" swimtime="00:00:35.90"/></SPLITS></RESULT><RESULT eventid="27" heatid="270" lane="1" points="434" resultid="2003" swimtime="00:00:35.62"><SPLITS/></RESULT><RESULT eventid="29" heatid="305" lane="1" points="454" resultid="2269" swimtime="00:02:26.98"><SPLITS><SPLIT distance="50" swimtime="00:00:32.60"/><SPLIT distance="100" swimtime="00:01:09.28"/><SPLIT distance="150" swimtime="00:01:48.01"/></SPLITS></RESULT><RESULT eventid="37" heatid="411" lane="1" points="478" resultid="3063" swimtime="00:02:37.70"><SPLITS><SPLIT distance="100" swimtime="00:01:16.87"/></SPLITS></RESULT><RESULT eventid="39" heatid="445" lane="6" points="457" resultid="3326" swimtime="00:01:07.10"><SPLITS><SPLIT distance="50" swimtime="00:00:31.90"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="382" birthdate="2014-01-01" firstname="Elias" gender="M" lastname="Klein" license="460784"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="54" lane="2" points="172" resultid="403" swimtime="00:06:35.33"><SPLITS><SPLIT distance="100" swimtime="00:01:33.08"/><SPLIT distance="200" swimtime="00:03:15.96"/><SPLIT distance="300" swimtime="00:04:58.46"/></SPLITS></RESULT><RESULT eventid="12" heatid="176" lane="4" points="168" resultid="1331" swimtime="00:03:26.20"><SPLITS><SPLIT distance="50" swimtime="00:00:49.58"/><SPLIT distance="100" swimtime="00:01:38.92"/><SPLIT distance="150" swimtime="00:02:42.48"/></SPLITS></RESULT><RESULT eventid="14" heatid="216" lane="3" points="165" resultid="1637" swimtime="00:01:33.91"><SPLITS/></RESULT><RESULT eventid="30" heatid="312" lane="1" points="177" resultid="2319" swimtime="00:03:01.37"><SPLITS><SPLIT distance="50" swimtime="00:00:40.56"/><SPLIT distance="100" swimtime="00:01:27.99"/><SPLIT distance="150" swimtime="00:02:16.28"/></SPLITS></RESULT><RESULT eventid="38" heatid="414" lane="3" points="185" resultid="3085" swimtime="00:03:16.38"><SPLITS><SPLIT distance="100" swimtime="00:01:36.89"/><SPLIT distance="150" swimtime="00:02:29.27"/></SPLITS></RESULT><RESULT eventid="40" heatid="458" lane="8" points="174" resultid="3428" swimtime="00:01:23.78"><SPLITS><SPLIT distance="50" swimtime="00:00:39.93"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="383" birthdate="2015-01-01" firstname="Keno" gender="M" lastname="von Szczytnicki" license="488396"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="54" lane="4" points="167" resultid="405" swimtime="00:06:38.95"><SPLITS><SPLIT distance="100" swimtime="00:01:32.06"/><SPLIT distance="200" swimtime="00:03:14.73"/><SPLIT distance="300" swimtime="00:04:57.99"/></SPLITS></RESULT><RESULT eventid="12" heatid="176" lane="5" points="155" resultid="1332" swimtime="00:03:32.12"><SPLITS><SPLIT distance="50" swimtime="00:00:49.47"/><SPLIT distance="100" swimtime="00:01:41.04"/><SPLIT distance="150" swimtime="00:02:44.87"/></SPLITS></RESULT><RESULT eventid="14" heatid="217" lane="2" points="139" resultid="1644" swimtime="00:01:39.59"><SPLITS><SPLIT distance="50" swimtime="00:00:48.30"/></SPLITS></RESULT><RESULT eventid="28" heatid="279" lane="4" points="154" resultid="2072" swimtime="00:00:44.14"><SPLITS/></RESULT><RESULT eventid="30" heatid="313" lane="7" points="159" resultid="2332" swimtime="00:03:08.09"><SPLITS><SPLIT distance="50" swimtime="00:00:43.10"/><SPLIT distance="100" swimtime="00:01:32.58"/><SPLIT distance="150" swimtime="00:02:21.05"/></SPLITS></RESULT><RESULT eventid="36" heatid="388" lane="2" points="123" resultid="2887" swimtime="00:00:44.68"><SPLITS/></RESULT><RESULT eventid="38" heatid="415" lane="7" points="172" resultid="3097" swimtime="00:03:20.91"><SPLITS><SPLIT distance="50" swimtime="00:00:46.85"/><SPLIT distance="100" swimtime="00:01:40.64"/><SPLIT distance="150" swimtime="00:02:32.58"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="386" birthdate="2015-01-01" firstname="Levi" gender="M" lastname="Hofweber" license="465153"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="54" lane="7" points="165" resultid="408" swimtime="00:06:40.83"><SPLITS><SPLIT distance="100" swimtime="00:01:33.15"/><SPLIT distance="200" swimtime="00:03:18.11"/><SPLIT distance="300" swimtime="00:05:01.15"/></SPLITS></RESULT><RESULT eventid="12" heatid="176" lane="2" points="135" resultid="1329" swimtime="00:03:42.18"><SPLITS><SPLIT distance="50" swimtime="00:00:56.60"/><SPLIT distance="100" swimtime="00:01:50.38"/><SPLIT distance="150" swimtime="00:02:54.45"/></SPLITS></RESULT><RESULT eventid="14" heatid="216" lane="8" points="133" resultid="1642" swimtime="00:01:40.94"><SPLITS><SPLIT distance="50" swimtime="00:00:49.93"/></SPLITS></RESULT><RESULT eventid="28" heatid="279" lane="1" points="149" resultid="2069" swimtime="00:00:44.69"><SPLITS/></RESULT><RESULT eventid="30" heatid="312" lane="7" points="142" resultid="2325" swimtime="00:03:15.21"><SPLITS><SPLIT distance="50" swimtime="00:00:44.71"/><SPLIT distance="100" swimtime="00:01:36.14"/><SPLIT distance="150" swimtime="00:02:27.12"/></SPLITS></RESULT><RESULT eventid="38" heatid="415" lane="2" points="157" resultid="3092" swimtime="00:03:27.45"><SPLITS><SPLIT distance="50" swimtime="00:00:49.59"/><SPLIT distance="100" swimtime="00:01:43.30"/><SPLIT distance="150" swimtime="00:02:37.37"/></SPLITS></RESULT><RESULT eventid="40" heatid="456" lane="2" points="144" resultid="3407" swimtime="00:01:29.40"><SPLITS><SPLIT distance="50" swimtime="00:00:43.28"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="396" birthdate="2011-01-01" firstname="Mads Christian" gender="M" lastname="Gutschmidt" license="424970"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="56" lane="3" resultid="420" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="10" heatid="142" lane="6" resultid="1072" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="14" heatid="219" lane="6" resultid="1664" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="28" heatid="281" lane="6" resultid="2090" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="30" heatid="316" lane="8" resultid="2357" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="38" heatid="417" lane="8" resultid="3113" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="40" heatid="461" lane="7" resultid="3450" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="398" birthdate="2011-01-01" firstname="Rian" gender="M" lastname="O'Connell" license="424971"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="56" lane="7" points="206" resultid="424" swimtime="00:06:12.55"><SPLITS><SPLIT distance="100" swimtime="00:01:21.50"/><SPLIT distance="200" swimtime="00:02:57.05"/><SPLIT distance="300" swimtime="00:04:37.65"/></SPLITS></RESULT><RESULT eventid="10" heatid="142" lane="4" points="307" resultid="1070" swimtime="00:00:30.97"><SPLITS/></RESULT><RESULT eventid="14" heatid="219" lane="5" points="245" resultid="1663" swimtime="00:01:22.42"><SPLITS><SPLIT distance="50" swimtime="00:00:39.28"/></SPLITS></RESULT><RESULT eventid="28" heatid="283" lane="6" points="250" resultid="2106" swimtime="00:00:37.63"><SPLITS/></RESULT><RESULT eventid="30" heatid="316" lane="7" points="222" resultid="2356" swimtime="00:02:48.35"><SPLITS><SPLIT distance="50" swimtime="00:00:34.70"/><SPLIT distance="100" swimtime="00:01:16.47"/><SPLIT distance="150" swimtime="00:02:02.23"/></SPLITS></RESULT><RESULT eventid="38" heatid="416" lane="2" points="243" resultid="3100" swimtime="00:02:59.35"><SPLITS><SPLIT distance="50" swimtime="00:00:40.59"/><SPLIT distance="100" swimtime="00:01:25.64"/><SPLIT distance="150" swimtime="00:02:13.79"/></SPLITS></RESULT><RESULT eventid="40" heatid="461" lane="2" points="291" resultid="3445" swimtime="00:01:10.71"><SPLITS><SPLIT distance="50" swimtime="00:00:32.79"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="399" birthdate="2013-01-01" firstname="Maximilian" gender="M" lastname="Lanz" license="465021"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="56" lane="8" points="192" resultid="425" swimtime="00:06:20.95"><SPLITS><SPLIT distance="100" swimtime="00:01:27.06"/><SPLIT distance="200" swimtime="00:03:04.52"/><SPLIT distance="300" swimtime="00:04:44.59"/></SPLITS></RESULT><RESULT eventid="10" heatid="139" lane="7" points="209" resultid="1050" swimtime="00:00:35.20"><SPLITS/></RESULT><RESULT eventid="14" heatid="218" lane="6" points="207" resultid="1656" swimtime="00:01:27.14"><SPLITS><SPLIT distance="50" swimtime="00:00:43.05"/></SPLITS></RESULT><RESULT eventid="30" heatid="314" lane="2" points="191" resultid="2335" swimtime="00:02:56.94"><SPLITS><SPLIT distance="50" swimtime="00:00:39.71"/><SPLIT distance="100" swimtime="00:01:27.27"/><SPLIT distance="150" swimtime="00:02:13.79"/></SPLITS></RESULT><RESULT eventid="38" heatid="414" lane="4" points="200" resultid="3086" swimtime="00:03:11.25"><SPLITS><SPLIT distance="50" swimtime="00:00:45.09"/><SPLIT distance="100" swimtime="00:01:35.35"/><SPLIT distance="150" swimtime="00:02:25.48"/></SPLITS></RESULT><RESULT comment="16:54 Start vor dem Startsignal" eventid="40" heatid="458" lane="5" resultid="3425" status="DSQ" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="411" birthdate="2012-01-01" firstname="Maximilian" gender="M" lastname="Hirsch" license="436074"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="58" lane="7" points="312" resultid="440" swimtime="00:05:24.41"><SPLITS><SPLIT distance="100" swimtime="00:01:17.41"/><SPLIT distance="200" swimtime="00:02:41.48"/><SPLIT distance="300" swimtime="00:04:04.56"/></SPLITS></RESULT><RESULT eventid="10" heatid="143" lane="3" points="276" resultid="1076" swimtime="00:00:32.09"><SPLITS/></RESULT><RESULT eventid="12" heatid="182" lane="7" points="279" resultid="1380" swimtime="00:02:54.31"><SPLITS><SPLIT distance="50" swimtime="00:00:39.58"/><SPLIT distance="100" swimtime="00:01:24.45"/><SPLIT distance="150" swimtime="00:02:15.16"/></SPLITS></RESULT><RESULT eventid="30" heatid="316" lane="3" points="297" resultid="2352" swimtime="00:02:32.85"><SPLITS><SPLIT distance="50" swimtime="00:00:35.61"/><SPLIT distance="100" swimtime="00:01:15.04"/><SPLIT distance="150" swimtime="00:01:55.71"/></SPLITS></RESULT><RESULT eventid="36" heatid="389" lane="6" points="210" resultid="2899" swimtime="00:00:37.44"><SPLITS/></RESULT><RESULT eventid="40" heatid="465" lane="3" points="307" resultid="3477" swimtime="00:01:09.39"><SPLITS><SPLIT distance="50" swimtime="00:00:33.78"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="439" birthdate="2014-01-01" firstname="Victoria Sophia" gender="F" lastname="Wiegartner" license="460791"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="5" heatid="63" lane="5" points="137" resultid="471" swimtime="00:01:47.47"><SPLITS><SPLIT distance="50" swimtime="00:00:48.59"/></SPLITS></RESULT><RESULT eventid="11" heatid="160" lane="4" points="215" resultid="1206" swimtime="00:03:30.41"><SPLITS><SPLIT distance="50" swimtime="00:00:47.69"/><SPLIT distance="100" swimtime="00:01:39.38"/><SPLIT distance="150" swimtime="00:02:41.39"/></SPLITS></RESULT><RESULT eventid="13" heatid="198" lane="8" points="202" resultid="1503" swimtime="00:01:37.87"><SPLITS><SPLIT distance="50" swimtime="00:00:48.27"/></SPLITS></RESULT><RESULT eventid="29" heatid="294" lane="8" points="229" resultid="2189" swimtime="00:03:04.47"><SPLITS><SPLIT distance="50" swimtime="00:00:42.95"/><SPLIT distance="100" swimtime="00:01:28.99"/><SPLIT distance="150" swimtime="00:02:19.46"/></SPLITS></RESULT><RESULT eventid="37" heatid="402" lane="3" points="217" resultid="2994" swimtime="00:03:25.11"><SPLITS><SPLIT distance="50" swimtime="00:00:47.92"/><SPLIT distance="100" swimtime="00:01:40.01"/><SPLIT distance="150" swimtime="00:02:34.09"/></SPLITS></RESULT><RESULT eventid="39" heatid="428" lane="3" points="197" resultid="3188" swimtime="00:01:28.84"><SPLITS><SPLIT distance="50" swimtime="00:00:42.73"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="448" birthdate="2012-01-01" firstname="Franziska" gender="F" lastname="Claßen" license="436075"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="5" heatid="66" lane="2" points="310" resultid="490" swimtime="00:01:21.92"><SPLITS><SPLIT distance="50" swimtime="00:00:36.96"/></SPLITS></RESULT><RESULT eventid="9" heatid="120" lane="5" points="461" resultid="908" swimtime="00:00:30.63"><SPLITS/></RESULT><RESULT eventid="11" heatid="168" lane="2" points="391" resultid="1268" swimtime="00:02:52.40"><SPLITS><SPLIT distance="50" swimtime="00:00:39.41"/><SPLIT distance="100" swimtime="00:01:22.56"/><SPLIT distance="150" swimtime="00:02:14.71"/></SPLITS></RESULT><RESULT eventid="27" heatid="265" lane="6" points="410" resultid="1969" swimtime="00:00:36.30"><SPLITS/></RESULT><RESULT eventid="29" heatid="301" lane="7" points="442" resultid="2243" swimtime="00:02:28.27"><SPLITS><SPLIT distance="50" swimtime="00:00:34.23"/><SPLIT distance="100" swimtime="00:01:12.54"/><SPLIT distance="150" swimtime="00:01:50.76"/></SPLITS></RESULT><RESULT eventid="35" heatid="372" lane="7" points="322" resultid="2773" swimtime="00:00:35.61"><SPLITS/></RESULT><RESULT eventid="39" heatid="440" lane="3" points="463" resultid="3283" swimtime="00:01:06.83"><SPLITS><SPLIT distance="50" swimtime="00:00:32.83"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="450" birthdate="2013-01-01" firstname="Luna Elisabeth" gender="F" lastname="Oettrich" license="441353"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="5" heatid="67" lane="1" points="275" resultid="497" swimtime="00:01:25.27"><SPLITS><SPLIT distance="50" swimtime="00:00:40.18"/></SPLITS></RESULT><RESULT eventid="11" heatid="167" lane="3" points="374" resultid="1261" swimtime="00:02:55.01"><SPLITS><SPLIT distance="50" swimtime="00:00:39.20"/><SPLIT distance="100" swimtime="00:01:21.75"/><SPLIT distance="150" swimtime="00:02:16.55"/></SPLITS></RESULT><RESULT eventid="13" heatid="202" lane="3" points="372" resultid="1530" swimtime="00:01:19.88"><SPLITS><SPLIT distance="50" swimtime="00:00:38.27"/></SPLITS></RESULT><RESULT eventid="27" heatid="265" lane="8" points="401" resultid="1971" swimtime="00:00:36.58"><SPLITS/></RESULT><RESULT eventid="37" heatid="407" lane="6" points="371" resultid="3036" swimtime="00:02:51.61"><SPLITS><SPLIT distance="50" swimtime="00:00:40.35"/><SPLIT distance="100" swimtime="00:01:24.68"/><SPLIT distance="150" swimtime="00:02:08.47"/></SPLITS></RESULT><RESULT eventid="39" heatid="438" lane="7" points="383" resultid="3272" swimtime="00:01:11.16"><SPLITS><SPLIT distance="50" swimtime="00:00:32.94"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="451" birthdate="2008-01-01" firstname="Carlotta" gender="F" lastname="Ambrosini" license="389645"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="5" heatid="67" lane="6" points="301" resultid="501" swimtime="00:01:22.74"><SPLITS><SPLIT distance="50" swimtime="00:00:37.22"/></SPLITS></RESULT><RESULT eventid="9" heatid="117" lane="5" points="408" resultid="884" swimtime="00:00:31.90"><SPLITS/></RESULT><RESULT eventid="13" heatid="206" lane="2" points="427" resultid="1561" swimtime="00:01:16.29"><SPLITS><SPLIT distance="50" swimtime="00:00:37.21"/></SPLITS></RESULT><RESULT eventid="27" heatid="268" lane="2" points="413" resultid="1989" swimtime="00:00:36.22"><SPLITS/></RESULT><RESULT eventid="35" heatid="375" lane="6" points="364" resultid="2795" swimtime="00:00:34.19"><SPLITS/></RESULT><RESULT eventid="37" heatid="410" lane="3" points="447" resultid="3057" swimtime="00:02:41.25"><SPLITS><SPLIT distance="50" swimtime="00:00:38.27"/><SPLIT distance="100" swimtime="00:01:18.65"/><SPLIT distance="150" swimtime="00:02:00.74"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="472" birthdate="2012-01-01" firstname="Alexander Silin" gender="M" lastname="Shen" license="436070"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="6" heatid="73" lane="2" points="253" resultid="545" swimtime="00:01:18.17"><SPLITS><SPLIT distance="50" swimtime="00:00:35.66"/></SPLITS></RESULT><RESULT eventid="10" heatid="144" lane="3" points="325" resultid="1084" swimtime="00:00:30.39"><SPLITS/></RESULT><RESULT eventid="12" heatid="183" lane="5" points="355" resultid="1386" swimtime="00:02:40.94"><SPLITS><SPLIT distance="50" swimtime="00:00:36.46"/><SPLIT distance="100" swimtime="00:01:18.44"/><SPLIT distance="150" swimtime="00:02:04.34"/></SPLITS></RESULT><RESULT eventid="28" heatid="282" lane="4" points="285" resultid="2096" swimtime="00:00:36.00"><SPLITS/></RESULT><RESULT eventid="30" heatid="319" lane="8" points="330" resultid="2381" swimtime="00:02:27.54"><SPLITS><SPLIT distance="50" swimtime="00:00:33.85"/><SPLIT distance="100" swimtime="00:01:11.77"/><SPLIT distance="150" swimtime="00:01:51.29"/></SPLITS></RESULT><RESULT eventid="36" heatid="390" lane="6" points="274" resultid="2907" swimtime="00:00:34.28"><SPLITS/></RESULT><RESULT eventid="40" heatid="465" lane="7" points="349" resultid="3481" swimtime="00:01:06.54"><SPLITS><SPLIT distance="50" swimtime="00:00:31.41"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="476" birthdate="2011-01-01" firstname="Anton" gender="M" lastname="Willmann" license="424964"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="6" heatid="73" lane="8" points="178" resultid="550" swimtime="00:01:27.88"><SPLITS><SPLIT distance="50" swimtime="00:00:40.39"/></SPLITS></RESULT><RESULT eventid="10" heatid="144" lane="7" points="331" resultid="1088" swimtime="00:00:30.22"><SPLITS/></RESULT><RESULT eventid="12" heatid="180" lane="6" points="269" resultid="1363" swimtime="00:02:56.57"><SPLITS><SPLIT distance="50" swimtime="00:00:38.84"/><SPLIT distance="100" swimtime="00:01:24.97"/><SPLIT distance="150" swimtime="00:02:18.49"/></SPLITS></RESULT><RESULT eventid="30" heatid="317" lane="6" points="259" resultid="2363" swimtime="00:02:39.91"><SPLITS><SPLIT distance="50" swimtime="00:00:35.03"/><SPLIT distance="100" swimtime="00:01:15.22"/><SPLIT distance="150" swimtime="00:01:59.10"/></SPLITS></RESULT><RESULT eventid="36" heatid="389" lane="2" points="236" resultid="2895" swimtime="00:00:35.99"><SPLITS/></RESULT><RESULT eventid="40" heatid="463" lane="4" points="325" resultid="3462" swimtime="00:01:08.14"><SPLITS><SPLIT distance="50" swimtime="00:00:32.27"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="485" birthdate="2009-01-01" firstname="Pascal" gender="M" lastname="van der Linden" license="411700"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="6" heatid="76" lane="4" points="352" resultid="570" swimtime="00:01:10.02"><SPLITS><SPLIT distance="50" swimtime="00:00:31.63"/></SPLITS></RESULT><RESULT eventid="10" heatid="150" lane="8" points="403" resultid="1137" swimtime="00:00:28.29"><SPLITS/></RESULT><RESULT eventid="14" heatid="224" lane="1" points="397" resultid="1697" swimtime="00:01:10.17"><SPLITS><SPLIT distance="50" swimtime="00:00:33.97"/></SPLITS></RESULT><RESULT eventid="28" heatid="285" lane="4" points="446" resultid="2119" swimtime="00:00:31.02"><SPLITS/></RESULT><RESULT eventid="36" heatid="394" lane="4" points="419" resultid="2937" swimtime="00:00:29.74"><SPLITS/></RESULT><RESULT eventid="38" heatid="419" lane="8" points="402" resultid="3126" swimtime="00:02:31.54"><SPLITS><SPLIT distance="50" swimtime="00:00:35.01"/><SPLIT distance="100" swimtime="00:01:13.09"/><SPLIT distance="150" swimtime="00:01:52.89"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="499" birthdate="2008-01-01" firstname="Jakob" gender="M" lastname="Seyfert" license="382545"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="6" heatid="79" lane="6" resultid="595" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="10" heatid="153" lane="3" resultid="1156" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="12" heatid="186" lane="4" resultid="1407" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="30" heatid="323" lane="8" resultid="2410" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="36" heatid="399" lane="8" resultid="2981" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="40" heatid="471" lane="2" resultid="3523" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="503" birthdate="1996-01-01" firstname="Dominik" gender="M" lastname="Liguori" license="180738"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="6" heatid="80" lane="6" points="569" resultid="602" swimtime="00:00:59.67"><SPLITS><SPLIT distance="50" swimtime="00:00:27.58"/></SPLITS></RESULT><RESULT eventid="10" heatid="157" lane="3" points="572" resultid="1186" swimtime="00:00:25.18"><SPLITS/></RESULT><RESULT eventid="12" heatid="189" lane="4" points="591" resultid="1431" swimtime="00:02:15.77"><SPLITS><SPLIT distance="50" swimtime="00:00:28.52"/><SPLIT distance="100" swimtime="00:01:05.06"/><SPLIT distance="150" swimtime="00:01:44.39"/></SPLITS></RESULT><RESULT eventid="30" heatid="325" lane="4" points="605" resultid="2421" swimtime="00:02:00.57"><SPLITS><SPLIT distance="50" swimtime="00:00:28.04"/><SPLIT distance="100" swimtime="00:00:58.90"/><SPLIT distance="150" swimtime="00:01:30.25"/></SPLITS></RESULT><RESULT eventid="36" heatid="400" lane="2" points="564" resultid="2982" swimtime="00:00:26.95"><SPLITS/></RESULT><RESULT eventid="40" heatid="475" lane="5" points="636" resultid="3556" swimtime="00:00:54.47"><SPLITS><SPLIT distance="50" swimtime="00:00:26.51"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="541" birthdate="2015-01-01" firstname="Valentin" gender="M" lastname="Li" license="465022"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="10" heatid="136" lane="8" points="93" resultid="1028" swimtime="00:00:46.05"><SPLITS/></RESULT><RESULT eventid="14" heatid="214" lane="3" points="139" resultid="1623" swimtime="00:01:39.40"><SPLITS><SPLIT distance="50" swimtime="00:00:48.21"/></SPLITS></RESULT><RESULT eventid="28" heatid="278" lane="8" points="107" resultid="2068" swimtime="00:00:49.79"><SPLITS/></RESULT><RESULT eventid="30" heatid="310" lane="1" points="116" resultid="2304" swimtime="00:03:28.72"><SPLITS><SPLIT distance="50" swimtime="00:00:48.10"/><SPLIT distance="100" swimtime="00:01:44.36"/><SPLIT distance="150" swimtime="00:02:39.51"/></SPLITS></RESULT><RESULT comment="15:31 Der Sportler hat bei der 100m Wende mehr als den einen erlaubten Armzug in Bauchlage ausgeführt" eventid="38" heatid="413" lane="6" resultid="3081" status="DSQ" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="40" heatid="454" lane="3" points="116" resultid="3392" swimtime="00:01:35.99"><SPLITS><SPLIT distance="50" swimtime="00:00:48.92"/></SPLITS></RESULT></RESULTS></ATHLETE></ATHLETES><RELAYS/></CLUB><CLUB code="4452" name="TSV Hohenbrunn-Riemerling" nation="GER" region="02" shortname="Hohenbrn" type="CLUB"><CONTACT city="Baiern" country="GER" email="kathi-schweiger@outlook.de" name="Schweiger, Katharina" phone="01522/9849011" street="Bergstraße 41" zip="85625"/><OFFICIALS/><ATHLETES><ATHLETE athleteid="32" birthdate="2015-01-01" firstname="Lynn" gender="F" lastname="Ossmann" license="466112"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="5" lane="4" points="172" resultid="32" swimtime="00:00:52.61"><SPLITS/></RESULT><RESULT eventid="7" heatid="81" lane="4" points="225" resultid="607" swimtime="00:03:48.33"><SPLITS><SPLIT distance="50" swimtime="00:00:54.88"/><SPLIT distance="100" swimtime="00:01:53.00"/><SPLIT distance="150" swimtime="00:02:51.46"/></SPLITS></RESULT><RESULT eventid="9" heatid="113" lane="5" points="288" resultid="853" swimtime="00:00:35.83"><SPLITS/></RESULT><RESULT eventid="13" heatid="197" lane="5" points="256" resultid="1492" swimtime="00:01:30.41"><SPLITS><SPLIT distance="50" swimtime="00:00:45.37"/></SPLITS></RESULT><RESULT eventid="27" heatid="261" lane="4" points="260" resultid="1935" swimtime="00:00:42.26"><SPLITS/></RESULT><RESULT eventid="31" heatid="329" lane="4" points="205" resultid="2446" swimtime="00:01:48.71"><SPLITS><SPLIT distance="50" swimtime="00:00:52.00"/></SPLITS></RESULT><RESULT eventid="35" heatid="366" lane="3" points="201" resultid="2721" swimtime="00:00:41.70"><SPLITS/></RESULT><RESULT eventid="37" heatid="404" lane="1" points="283" resultid="3007" swimtime="00:03:07.79"><SPLITS><SPLIT distance="50" swimtime="00:00:46.58"/><SPLIT distance="100" swimtime="00:01:34.24"/><SPLIT distance="150" swimtime="00:02:23.88"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="37" birthdate="2015-01-01" firstname="Inessa" gender="F" lastname="Elbing" license="483053"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="6" lane="1" points="142" resultid="37" swimtime="00:00:56.12"><SPLITS/></RESULT><RESULT eventid="9" heatid="109" lane="5" points="196" resultid="821" swimtime="00:00:40.71"><SPLITS/></RESULT><RESULT eventid="11" heatid="158" lane="4" points="177" resultid="1193" swimtime="00:03:44.49"><SPLITS><SPLIT distance="50" swimtime="00:00:51.76"/><SPLIT distance="100" swimtime="00:01:49.06"/><SPLIT distance="150" swimtime="00:02:56.07"/></SPLITS></RESULT><RESULT eventid="29" heatid="291" lane="8" points="200" resultid="2165" swimtime="00:03:13.16"><SPLITS><SPLIT distance="50" swimtime="00:00:44.02"/><SPLIT distance="100" swimtime="00:01:32.69"/><SPLIT distance="150" swimtime="00:02:26.24"/></SPLITS></RESULT><RESULT eventid="35" heatid="364" lane="8" points="107" resultid="2710" swimtime="00:00:51.43"><SPLITS/></RESULT><RESULT eventid="37" heatid="402" lane="5" points="162" resultid="2996" swimtime="00:03:46.05"><SPLITS><SPLIT distance="50" swimtime="00:00:54.32"/><SPLIT distance="100" swimtime="00:01:54.23"/></SPLITS></RESULT><RESULT eventid="39" heatid="427" lane="7" points="176" resultid="3184" swimtime="00:01:32.25"><SPLITS><SPLIT distance="50" swimtime="00:00:44.51"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="53" birthdate="2014-01-01" firstname="Anouk" gender="F" lastname="Stevenson" license="490223"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="8" lane="1" points="178" resultid="53" swimtime="00:00:52.07"><SPLITS/></RESULT><RESULT eventid="7" heatid="81" lane="3" points="206" resultid="606" swimtime="00:03:55.01"><SPLITS><SPLIT distance="50" swimtime="00:00:54.06"/><SPLIT distance="100" swimtime="00:01:54.47"/><SPLIT distance="150" swimtime="00:02:56.89"/></SPLITS></RESULT><RESULT eventid="9" heatid="107" lane="6" points="161" resultid="806" swimtime="00:00:43.44"><SPLITS/></RESULT><RESULT eventid="13" heatid="191" lane="1" points="127" resultid="1440" swimtime="00:01:54.10"><SPLITS><SPLIT distance="50" swimtime="00:00:56.92"/></SPLITS></RESULT><RESULT eventid="23" heatid="241" lane="7" resultid="1798" swimtime="00:01:13.72"><SPLITS/></RESULT><RESULT eventid="25" heatid="247" lane="5" resultid="1834" swimtime="00:01:02.80"><SPLITS/></RESULT><RESULT eventid="31" heatid="330" lane="1" points="176" resultid="2451" swimtime="00:01:54.34"><SPLITS/></RESULT><RESULT eventid="39" heatid="423" lane="6" points="127" resultid="3152" swimtime="00:01:42.61"><SPLITS><SPLIT distance="50" swimtime="00:00:47.74"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="55" birthdate="2014-01-01" firstname="Alma" gender="F" lastname="Scheithauer" license="483085"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="8" lane="3" points="186" resultid="55" swimtime="00:00:51.30"><SPLITS/></RESULT><RESULT eventid="7" heatid="84" lane="6" points="207" resultid="630" swimtime="00:03:54.88"><SPLITS><SPLIT distance="50" swimtime="00:00:49.90"/><SPLIT distance="100" swimtime="00:01:50.03"/><SPLIT distance="150" swimtime="00:02:51.81"/></SPLITS></RESULT><RESULT eventid="9" heatid="107" lane="5" points="164" resultid="805" swimtime="00:00:43.20"><SPLITS/></RESULT><RESULT eventid="13" heatid="190" lane="4" points="109" resultid="1437" swimtime="00:01:59.97"><SPLITS><SPLIT distance="50" swimtime="00:00:56.20"/></SPLITS></RESULT><RESULT eventid="19" heatid="234" lane="3" resultid="1759" swimtime="00:01:19.40"><SPLITS/></RESULT><RESULT eventid="25" heatid="247" lane="4" resultid="1833" swimtime="00:01:01.43"><SPLITS/></RESULT><RESULT eventid="31" heatid="333" lane="3" points="182" resultid="2477" swimtime="00:01:53.00"><SPLITS><SPLIT distance="50" swimtime="00:00:54.38"/></SPLITS></RESULT><RESULT eventid="39" heatid="421" lane="4" points="113" resultid="3134" swimtime="00:01:46.85"><SPLITS><SPLIT distance="50" swimtime="00:00:47.83"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="59" birthdate="2014-01-01" firstname="Rebekka" gender="F" lastname="Holland" license="483062"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="8" lane="7" points="167" resultid="59" swimtime="00:00:53.20"><SPLITS/></RESULT><RESULT eventid="7" heatid="81" lane="5" points="173" resultid="608" swimtime="00:04:08.99"><SPLITS><SPLIT distance="50" swimtime="00:00:56.38"/><SPLIT distance="100" swimtime="00:02:00.81"/><SPLIT distance="150" swimtime="00:03:05.81"/></SPLITS></RESULT><RESULT eventid="9" heatid="108" lane="8" points="133" resultid="816" swimtime="00:00:46.35"><SPLITS/></RESULT><RESULT eventid="13" heatid="194" lane="1" points="147" resultid="1464" swimtime="00:01:48.62"><SPLITS><SPLIT distance="50" swimtime="00:00:54.30"/></SPLITS></RESULT><RESULT eventid="23" heatid="242" lane="5" resultid="1803" swimtime="00:01:02.28"><SPLITS/></RESULT><RESULT eventid="25" heatid="248" lane="8" resultid="1844" swimtime="00:01:05.28"><SPLITS/></RESULT><RESULT eventid="29" heatid="289" lane="7" points="107" resultid="2149" swimtime="00:03:57.33"><SPLITS><SPLIT distance="50" swimtime="00:00:50.51"/><SPLIT distance="100" swimtime="00:01:53.27"/><SPLIT distance="150" swimtime="00:02:57.12"/></SPLITS></RESULT><RESULT eventid="35" heatid="364" lane="5" points="82" resultid="2707" swimtime="00:00:56.20"><SPLITS/></RESULT><RESULT eventid="39" heatid="423" lane="2" points="100" resultid="3148" swimtime="00:01:51.08"><SPLITS><SPLIT distance="50" swimtime="00:00:51.34"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="66" birthdate="2013-01-01" firstname="Theresa" gender="F" lastname="Schramm" license="490081"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="9" lane="6" points="206" resultid="66" swimtime="00:00:49.56"><SPLITS/></RESULT><RESULT eventid="7" heatid="81" lane="6" points="193" resultid="609" swimtime="00:04:00.35"><SPLITS><SPLIT distance="50" swimtime="00:00:54.85"/><SPLIT distance="100" swimtime="00:01:57.42"/><SPLIT distance="150" swimtime="00:03:01.59"/></SPLITS></RESULT><RESULT eventid="9" heatid="109" lane="7" points="195" resultid="823" swimtime="00:00:40.77"><SPLITS/></RESULT><RESULT eventid="13" heatid="193" lane="6" points="140" resultid="1461" swimtime="00:01:50.55"><SPLITS><SPLIT distance="50" swimtime="00:00:52.30"/></SPLITS></RESULT><RESULT eventid="23" heatid="240" lane="4" resultid="1791" swimtime="00:01:01.74"><SPLITS/></RESULT><RESULT eventid="25" heatid="247" lane="3" resultid="1832" swimtime="00:01:00.52"><SPLITS/></RESULT><RESULT eventid="31" heatid="332" lane="7" points="191" resultid="2473" swimtime="00:01:51.27"><SPLITS><SPLIT distance="50" swimtime="00:00:52.63"/></SPLITS></RESULT><RESULT eventid="39" heatid="425" lane="4" points="149" resultid="3166" swimtime="00:01:37.45"><SPLITS><SPLIT distance="50" swimtime="00:00:45.70"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="86" birthdate="2015-01-01" firstname="Azzurra" gender="F" lastname="Dostetan Affuso" license="464843"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="12" lane="2" points="178" resultid="86" swimtime="00:00:52.00"><SPLITS/></RESULT><RESULT eventid="7" heatid="84" lane="8" points="174" resultid="632" swimtime="00:04:08.79"><SPLITS><SPLIT distance="50" swimtime="00:00:58.78"/><SPLIT distance="100" swimtime="00:02:00.20"/><SPLIT distance="150" swimtime="00:03:09.89"/></SPLITS></RESULT><RESULT eventid="9" heatid="110" lane="5" points="196" resultid="829" swimtime="00:00:40.73"><SPLITS/></RESULT><RESULT eventid="11" heatid="158" lane="5" points="168" resultid="1194" swimtime="00:03:48.35"><SPLITS><SPLIT distance="50" swimtime="00:00:57.39"/><SPLIT distance="100" swimtime="00:01:53.87"/><SPLIT distance="150" swimtime="00:02:59.02"/></SPLITS></RESULT><RESULT eventid="29" heatid="291" lane="6" points="180" resultid="2163" swimtime="00:03:20.06"><SPLITS><SPLIT distance="50" swimtime="00:00:44.37"/><SPLIT distance="100" swimtime="00:01:36.64"/><SPLIT distance="150" swimtime="00:02:30.65"/></SPLITS></RESULT><RESULT eventid="31" heatid="330" lane="5" points="162" resultid="2455" swimtime="00:01:57.54"><SPLITS/></RESULT><RESULT eventid="35" heatid="365" lane="8" points="84" resultid="2718" swimtime="00:00:55.72"><SPLITS/></RESULT><RESULT eventid="39" heatid="429" lane="8" points="177" resultid="3201" swimtime="00:01:31.98"><SPLITS><SPLIT distance="50" swimtime="00:00:43.91"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="87" birthdate="2014-01-01" firstname="Sophia" gender="F" lastname="Wild" license="483747"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="12" lane="3" resultid="87" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="7" heatid="84" lane="4" resultid="628" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="9" heatid="109" lane="2" resultid="818" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="13" heatid="193" lane="7" resultid="1462" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="23" heatid="242" lane="3" resultid="1801" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="25" heatid="249" lane="8" resultid="1852" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="31" heatid="334" lane="3" resultid="2485" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="35" heatid="363" lane="4" resultid="2698" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="92" birthdate="2013-01-01" firstname="Katharina" gender="F" lastname="Lang" license="483068"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="12" lane="8" points="229" resultid="92" swimtime="00:00:47.83"><SPLITS/></RESULT><RESULT eventid="7" heatid="85" lane="7" points="267" resultid="639" swimtime="00:03:35.71"><SPLITS><SPLIT distance="50" swimtime="00:00:49.21"/><SPLIT distance="100" swimtime="00:01:45.35"/><SPLIT distance="150" swimtime="00:02:41.15"/></SPLITS></RESULT><RESULT eventid="11" heatid="161" lane="4" points="260" resultid="1214" swimtime="00:03:17.59"><SPLITS><SPLIT distance="50" swimtime="00:00:43.09"/><SPLIT distance="100" swimtime="00:01:34.14"/><SPLIT distance="150" swimtime="00:02:30.26"/></SPLITS></RESULT><RESULT eventid="13" heatid="199" lane="3" points="232" resultid="1506" swimtime="00:01:33.47"><SPLITS><SPLIT distance="50" swimtime="00:00:46.91"/></SPLITS></RESULT><RESULT eventid="19" heatid="234" lane="4" resultid="1760" swimtime="00:01:02.10"><SPLITS/></RESULT><RESULT eventid="27" heatid="261" lane="7" points="241" resultid="1938" swimtime="00:00:43.31"><SPLITS/></RESULT><RESULT eventid="31" heatid="334" lane="8" points="250" resultid="2490" swimtime="00:01:41.80"><SPLITS><SPLIT distance="50" swimtime="00:00:49.40"/></SPLITS></RESULT><RESULT eventid="35" heatid="367" lane="3" points="160" resultid="2729" swimtime="00:00:44.97"><SPLITS/></RESULT><RESULT eventid="37" heatid="405" lane="5" resultid="3019" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="103" birthdate="2013-01-01" firstname="Hannah" gender="F" lastname="Janosek" license="483066"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="14" lane="3" points="252" resultid="103" swimtime="00:00:46.38"><SPLITS/></RESULT><RESULT eventid="5" heatid="64" lane="5" points="199" resultid="477" swimtime="00:01:34.88"><SPLITS><SPLIT distance="50" swimtime="00:00:43.74"/></SPLITS></RESULT><RESULT eventid="11" heatid="165" lane="8" points="276" resultid="1250" swimtime="00:03:13.63"><SPLITS><SPLIT distance="50" swimtime="00:00:43.41"/><SPLIT distance="100" swimtime="00:01:32.08"/><SPLIT distance="150" swimtime="00:02:31.58"/></SPLITS></RESULT><RESULT eventid="13" heatid="201" lane="8" points="260" resultid="1527" swimtime="00:01:29.98"><SPLITS><SPLIT distance="50" swimtime="00:00:42.79"/></SPLITS></RESULT><RESULT eventid="21" heatid="238" lane="7" resultid="1784" swimtime="00:01:05.41"><SPLITS/></RESULT><RESULT eventid="27" heatid="262" lane="3" points="295" resultid="1942" swimtime="00:00:40.49"><SPLITS/></RESULT><RESULT eventid="31" heatid="336" lane="4" points="243" resultid="2502" swimtime="00:01:42.72"><SPLITS><SPLIT distance="50" swimtime="00:00:47.69"/></SPLITS></RESULT><RESULT eventid="35" heatid="369" lane="4" points="237" resultid="2746" swimtime="00:00:39.47"><SPLITS/></RESULT><RESULT eventid="37" heatid="406" lane="7" points="274" resultid="3029" swimtime="00:03:09.74"><SPLITS><SPLIT distance="50" swimtime="00:00:44.17"/><SPLIT distance="100" swimtime="00:01:33.48"/><SPLIT distance="150" swimtime="00:02:22.72"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="112" birthdate="2014-01-01" firstname="Charlotte" gender="F" lastname="Schneider" license="490161"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="15" lane="4" points="274" resultid="112" swimtime="00:00:45.09"><SPLITS/></RESULT><RESULT eventid="9" heatid="115" lane="3" points="269" resultid="867" swimtime="00:00:36.65"><SPLITS/></RESULT><RESULT eventid="11" heatid="161" lane="7" points="226" resultid="1217" swimtime="00:03:26.92"><SPLITS><SPLIT distance="50" swimtime="00:00:45.97"/><SPLIT distance="100" swimtime="00:01:40.74"/><SPLIT distance="150" swimtime="00:02:41.76"/></SPLITS></RESULT><RESULT eventid="13" heatid="197" lane="6" points="227" resultid="1493" swimtime="00:01:34.12"><SPLITS><SPLIT distance="50" swimtime="00:00:44.95"/></SPLITS></RESULT><RESULT eventid="23" heatid="243" lane="7" resultid="1813" swimtime="00:00:51.00"><SPLITS/></RESULT><RESULT eventid="25" heatid="248" lane="1" resultid="1837" swimtime="00:01:00.70"><SPLITS/></RESULT><RESULT eventid="31" heatid="335" lane="8" points="261" resultid="2498" swimtime="00:01:40.27"><SPLITS><SPLIT distance="50" swimtime="00:00:48.87"/></SPLITS></RESULT><RESULT eventid="35" heatid="365" lane="2" points="162" resultid="2712" swimtime="00:00:44.75"><SPLITS/></RESULT><RESULT eventid="39" heatid="431" lane="7" points="231" resultid="3216" swimtime="00:01:24.26"><SPLITS><SPLIT distance="50" swimtime="00:00:39.58"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="114" birthdate="2013-01-01" firstname="Yana Katharina" gender="F" lastname="Deixler" license="462723"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="15" lane="6" points="345" resultid="114" swimtime="00:00:41.74"><SPLITS/></RESULT><RESULT eventid="7" heatid="87" lane="7" points="333" resultid="655" swimtime="00:03:20.44"><SPLITS><SPLIT distance="50" swimtime="00:00:44.36"/><SPLIT distance="100" swimtime="00:01:35.25"/><SPLIT distance="150" swimtime="00:02:28.51"/></SPLITS></RESULT><RESULT eventid="9" heatid="113" lane="3" points="346" resultid="851" swimtime="00:00:33.69"><SPLITS/></RESULT><RESULT eventid="25" heatid="249" lane="2" resultid="1846" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="31" heatid="336" lane="5" points="336" resultid="2503" swimtime="00:01:32.23"><SPLITS><SPLIT distance="50" swimtime="00:00:43.53"/></SPLITS></RESULT><RESULT eventid="35" heatid="367" lane="7" resultid="2733" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="39" heatid="433" lane="3" points="329" resultid="3228" swimtime="00:01:14.86"><SPLITS><SPLIT distance="50" swimtime="00:00:35.98"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="116" birthdate="2014-01-01" firstname="Linnea" gender="F" lastname="Johnsson" license="483075"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="15" lane="8" points="231" resultid="116" swimtime="00:00:47.72"><SPLITS/></RESULT><RESULT eventid="7" heatid="86" lane="5" points="261" resultid="645" swimtime="00:03:37.28"><SPLITS><SPLIT distance="50" swimtime="00:00:46.99"/><SPLIT distance="100" swimtime="00:01:43.11"/><SPLIT distance="150" swimtime="00:02:40.79"/></SPLITS></RESULT><RESULT eventid="9" heatid="112" lane="1" points="231" resultid="841" swimtime="00:00:38.56"><SPLITS/></RESULT><RESULT eventid="13" heatid="199" lane="7" points="211" resultid="1510" swimtime="00:01:36.41"><SPLITS><SPLIT distance="50" swimtime="00:00:46.49"/></SPLITS></RESULT><RESULT eventid="23" heatid="243" lane="2" resultid="1808" swimtime="00:00:48.64"><SPLITS/></RESULT><RESULT eventid="25" heatid="249" lane="6" resultid="1850" swimtime="00:00:58.86"><SPLITS/></RESULT><RESULT eventid="31" heatid="335" lane="2" points="238" resultid="2492" swimtime="00:01:43.43"><SPLITS><SPLIT distance="50" swimtime="00:00:49.55"/></SPLITS></RESULT><RESULT eventid="35" heatid="365" lane="7" points="126" resultid="2717" swimtime="00:00:48.62"><SPLITS/></RESULT><RESULT eventid="37" heatid="404" lane="4" points="210" resultid="3010" swimtime="00:03:27.47"><SPLITS><SPLIT distance="50" swimtime="00:00:47.41"/><SPLIT distance="100" swimtime="00:01:42.03"/><SPLIT distance="150" swimtime="00:02:35.85"/></SPLITS></RESULT><RESULT eventid="39" heatid="428" lane="4" points="226" resultid="3189" swimtime="00:01:24.89"><SPLITS><SPLIT distance="50" swimtime="00:00:38.77"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="130" birthdate="2013-01-01" firstname="Zona" gender="F" lastname="Todorovic" license="483751"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="17" lane="6" points="364" resultid="130" swimtime="00:00:41.01"><SPLITS/></RESULT><RESULT eventid="7" heatid="88" lane="2" points="332" resultid="658" swimtime="00:03:20.51"><SPLITS><SPLIT distance="50" swimtime="00:00:44.25"/><SPLIT distance="100" swimtime="00:01:36.55"/><SPLIT distance="150" swimtime="00:02:30.90"/></SPLITS></RESULT><RESULT eventid="11" heatid="164" lane="1" points="285" resultid="1235" swimtime="00:03:11.60"><SPLITS><SPLIT distance="50" swimtime="00:00:45.98"/><SPLIT distance="100" swimtime="00:01:03.08"/><SPLIT distance="150" swimtime="00:02:32.10"/></SPLITS></RESULT><RESULT eventid="13" heatid="200" lane="1" points="268" resultid="1512" swimtime="00:01:29.10"><SPLITS><SPLIT distance="50" swimtime="00:00:43.72"/></SPLITS></RESULT><RESULT eventid="25" heatid="249" lane="1" resultid="1845" swimtime="00:00:57.75"><SPLITS/></RESULT><RESULT eventid="29" heatid="296" lane="3" points="325" resultid="2200" swimtime="00:02:44.22"><SPLITS><SPLIT distance="50" swimtime="00:00:37.80"/><SPLIT distance="100" swimtime="00:01:18.93"/><SPLIT distance="150" swimtime="00:02:02.67"/></SPLITS></RESULT><RESULT eventid="31" heatid="337" lane="3" points="327" resultid="2509" swimtime="00:01:33.04"><SPLITS><SPLIT distance="50" swimtime="00:00:44.63"/></SPLITS></RESULT><RESULT eventid="35" heatid="368" lane="8" points="153" resultid="2742" swimtime="00:00:45.59"><SPLITS/></RESULT><RESULT eventid="39" heatid="433" lane="5" points="339" resultid="3230" swimtime="00:01:14.13"><SPLITS><SPLIT distance="50" swimtime="00:00:36.18"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="171" birthdate="2011-01-01" firstname="Pia" gender="F" lastname="Junge" license="406943"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="23" lane="1" points="471" resultid="171" swimtime="00:00:37.65"><SPLITS/></RESULT><RESULT eventid="7" heatid="91" lane="8" points="464" resultid="688" swimtime="00:02:59.43"><SPLITS><SPLIT distance="50" swimtime="00:00:41.89"/><SPLIT distance="100" swimtime="00:01:28.33"/><SPLIT distance="150" swimtime="00:02:15.40"/></SPLITS></RESULT><RESULT eventid="9" heatid="123" lane="3" points="468" resultid="930" swimtime="00:00:30.48"><SPLITS/></RESULT><RESULT eventid="13" heatid="206" lane="3" points="440" resultid="1562" swimtime="00:01:15.53"><SPLITS><SPLIT distance="50" swimtime="00:00:36.90"/></SPLITS></RESULT><RESULT eventid="27" heatid="270" lane="2" points="500" resultid="2004" swimtime="00:00:33.99"><SPLITS/></RESULT><RESULT eventid="31" heatid="342" lane="2" points="451" resultid="2548" swimtime="00:01:23.62"><SPLITS><SPLIT distance="50" swimtime="00:00:39.52"/></SPLITS></RESULT><RESULT eventid="37" heatid="409" lane="7" points="439" resultid="3053" swimtime="00:02:42.19"><SPLITS><SPLIT distance="50" swimtime="00:00:37.92"/><SPLIT distance="100" swimtime="00:01:20.17"/><SPLIT distance="150" swimtime="00:02:02.39"/></SPLITS></RESULT><RESULT eventid="39" heatid="443" lane="3" points="438" resultid="3307" swimtime="00:01:08.07"><SPLITS><SPLIT distance="50" swimtime="00:00:32.75"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="181" birthdate="2011-01-01" firstname="Sophia" gender="F" lastname="Hofmann" license="406942"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="24" lane="3" points="436" resultid="181" swimtime="00:00:38.63"><SPLITS/></RESULT><RESULT eventid="5" heatid="69" lane="6" points="365" resultid="517" swimtime="00:01:17.61"><SPLITS><SPLIT distance="50" swimtime="00:00:34.81"/></SPLITS></RESULT><RESULT eventid="7" heatid="90" lane="2" points="446" resultid="674" swimtime="00:03:01.83"><SPLITS><SPLIT distance="50" swimtime="00:00:41.83"/><SPLIT distance="100" swimtime="00:01:27.91"/><SPLIT distance="150" swimtime="00:02:16.32"/></SPLITS></RESULT><RESULT eventid="9" heatid="128" lane="4" points="440" resultid="970" swimtime="00:00:31.12"><SPLITS/></RESULT><RESULT eventid="11" heatid="170" lane="5" points="413" resultid="1287" swimtime="00:02:49.28"><SPLITS><SPLIT distance="50" swimtime="00:00:35.44"/><SPLIT distance="100" swimtime="00:01:21.61"/><SPLIT distance="150" swimtime="00:02:10.01"/></SPLITS></RESULT><RESULT eventid="31" heatid="344" lane="2" points="465" resultid="2564" swimtime="00:01:22.76"><SPLITS><SPLIT distance="50" swimtime="00:00:38.76"/></SPLITS></RESULT><RESULT eventid="35" heatid="381" lane="5" points="392" resultid="2840" swimtime="00:00:33.38"><SPLITS/></RESULT><RESULT eventid="39" heatid="445" lane="3" points="445" resultid="3323" swimtime="00:01:07.73"><SPLITS><SPLIT distance="50" swimtime="00:00:32.86"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="183" birthdate="2010-01-01" firstname="Laura" gender="F" lastname="Gülzow" license="392671"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="24" lane="5" points="533" resultid="183" swimtime="00:00:36.13"><SPLITS/></RESULT><RESULT eventid="5" heatid="69" lane="5" points="408" resultid="516" swimtime="00:01:14.79"><SPLITS><SPLIT distance="50" swimtime="00:00:34.09"/></SPLITS></RESULT><RESULT eventid="7" heatid="91" lane="7" points="453" resultid="687" swimtime="00:03:00.81"><SPLITS><SPLIT distance="50" swimtime="00:00:42.13"/><SPLIT distance="100" swimtime="00:01:27.40"/><SPLIT distance="150" swimtime="00:02:13.45"/></SPLITS></RESULT><RESULT eventid="9" heatid="129" lane="1" points="450" resultid="975" swimtime="00:00:30.88"><SPLITS/></RESULT><RESULT eventid="11" heatid="171" lane="8" points="438" resultid="1298" swimtime="00:02:45.98"><SPLITS><SPLIT distance="50" swimtime="00:00:34.83"/><SPLIT distance="100" swimtime="00:01:21.69"/><SPLIT distance="150" swimtime="00:02:08.13"/></SPLITS></RESULT><RESULT eventid="31" heatid="344" lane="3" points="504" resultid="2565" swimtime="00:01:20.56"><SPLITS><SPLIT distance="50" swimtime="00:00:37.98"/></SPLITS></RESULT><RESULT eventid="35" heatid="380" lane="6" points="415" resultid="2833" swimtime="00:00:32.74"><SPLITS/></RESULT><RESULT eventid="39" heatid="448" lane="3" points="464" resultid="3345" swimtime="00:01:06.75"><SPLITS><SPLIT distance="50" swimtime="00:00:32.16"/></SPLITS></RESULT><RESULT eventid="41" heatid="477" lane="2" points="423" resultid="3564" swimtime="00:05:54.72"><SPLITS><SPLIT distance="50" swimtime="00:00:37.41"/><SPLIT distance="100" swimtime="00:01:20.86"/><SPLIT distance="150" swimtime="00:02:10.26"/><SPLIT distance="200" swimtime="00:02:58.31"/><SPLIT distance="250" swimtime="00:03:46.45"/><SPLIT distance="300" swimtime="00:04:33.34"/><SPLIT distance="350" swimtime="00:05:15.24"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="222" birthdate="2014-01-01" firstname="Jasper" gender="M" lastname="Nierbauer" license="483080"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="30" lane="2" points="105" resultid="222" swimtime="00:00:54.97"><SPLITS/></RESULT><RESULT eventid="8" heatid="94" lane="2" points="123" resultid="705" swimtime="00:04:12.97"><SPLITS><SPLIT distance="50" swimtime="00:00:57.14"/><SPLIT distance="100" swimtime="00:02:01.39"/><SPLIT distance="150" swimtime="00:03:07.58"/></SPLITS></RESULT><RESULT eventid="10" heatid="139" lane="6" points="160" resultid="1049" swimtime="00:00:38.46"><SPLITS/></RESULT><RESULT eventid="14" heatid="216" lane="7" points="142" resultid="1641" swimtime="00:01:38.74"><SPLITS><SPLIT distance="50" swimtime="00:00:46.61"/></SPLITS></RESULT><RESULT eventid="20" heatid="236" lane="2" resultid="1770" swimtime="00:01:07.65"><SPLITS/></RESULT><RESULT eventid="24" heatid="244" lane="5" resultid="1818" swimtime="00:01:05.09"><SPLITS/></RESULT><RESULT eventid="38" heatid="413" lane="2" points="165" resultid="3078" swimtime="00:03:23.85"><SPLITS><SPLIT distance="50" swimtime="00:00:49.03"/><SPLIT distance="100" swimtime="00:01:40.90"/><SPLIT distance="150" swimtime="00:02:35.22"/></SPLITS></RESULT><RESULT eventid="40" heatid="457" lane="8" points="137" resultid="3420" swimtime="00:01:30.84"><SPLITS><SPLIT distance="50" swimtime="00:00:41.95"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="223" birthdate="2015-01-01" firstname="Leo" gender="M" lastname="Alting van Geusau" license="483256"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="30" lane="3" points="123" resultid="223" swimtime="00:00:52.06"><SPLITS/></RESULT><RESULT eventid="8" heatid="96" lane="8" points="184" resultid="725" swimtime="00:03:41.26"><SPLITS><SPLIT distance="50" swimtime="00:00:51.95"/><SPLIT distance="100" swimtime="00:01:47.86"/><SPLIT distance="150" swimtime="00:02:45.59"/></SPLITS></RESULT><RESULT eventid="10" heatid="136" lane="7" points="132" resultid="1027" swimtime="00:00:40.99"><SPLITS/></RESULT><RESULT eventid="14" heatid="213" lane="6" points="122" resultid="1618" swimtime="00:01:43.77"><SPLITS><SPLIT distance="50" swimtime="00:00:50.17"/></SPLITS></RESULT><RESULT eventid="32" heatid="348" lane="1" points="145" resultid="2590" swimtime="00:01:48.15"><SPLITS><SPLIT distance="50" swimtime="00:00:53.70"/></SPLITS></RESULT><RESULT eventid="38" heatid="413" lane="5" resultid="3080" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="40" heatid="455" lane="1" points="139" resultid="3398" swimtime="00:01:30.43"><SPLITS><SPLIT distance="50" swimtime="00:00:43.15"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="225" birthdate="2014-01-01" firstname="Emil" gender="M" lastname="Seiler" license="483738"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="30" lane="5" points="128" resultid="225" swimtime="00:00:51.44"><SPLITS/></RESULT><RESULT eventid="8" heatid="93" lane="7" points="159" resultid="703" swimtime="00:03:52.05"><SPLITS><SPLIT distance="50" swimtime="00:00:52.62"/><SPLIT distance="100" swimtime="00:01:53.40"/><SPLIT distance="150" swimtime="00:02:54.77"/></SPLITS></RESULT><RESULT eventid="10" heatid="137" lane="3" points="152" resultid="1031" swimtime="00:00:39.10"><SPLITS/></RESULT><RESULT eventid="14" heatid="214" lane="5" points="138" resultid="1625" swimtime="00:01:39.68"><SPLITS><SPLIT distance="50" swimtime="00:00:49.13"/></SPLITS></RESULT><RESULT eventid="24" heatid="244" lane="6" resultid="1819" swimtime="00:00:56.13"><SPLITS/></RESULT><RESULT eventid="26" heatid="250" lane="4" resultid="1854" swimtime="00:01:01.18"><SPLITS/></RESULT><RESULT eventid="32" heatid="348" lane="2" points="124" resultid="2591" swimtime="00:01:53.92"><SPLITS><SPLIT distance="50" swimtime="00:00:56.78"/></SPLITS></RESULT><RESULT comment="14:27 Der Sportler führte mehrere Wechselbeinschläge aus" eventid="36" heatid="384" lane="2" resultid="2856" status="DSQ" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="40" heatid="455" lane="5" points="121" resultid="3402" swimtime="00:01:34.69"><SPLITS><SPLIT distance="50" swimtime="00:00:44.72"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="232" birthdate="2014-01-01" firstname="Björn" gender="M" lastname="Fuchs" license="477352"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="31" lane="4" points="166" resultid="232" swimtime="00:00:47.19"><SPLITS/></RESULT><RESULT eventid="6" heatid="72" lane="3" points="129" resultid="538" swimtime="00:01:37.62"><SPLITS><SPLIT distance="50" swimtime="00:00:44.79"/></SPLITS></RESULT><RESULT comment="16:13 Der Sportler hat beim Zielanschlag der Teilstrecke Schmetterling nicht mit beiden Händen gleichzeitig angeschlagen" eventid="12" heatid="178" lane="7" resultid="1348" status="DSQ" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="14" heatid="215" lane="7" points="152" resultid="1633" swimtime="00:01:36.58"><SPLITS><SPLIT distance="50" swimtime="00:00:47.03"/></SPLITS></RESULT><RESULT eventid="22" heatid="239" lane="6" resultid="1789" swimtime="00:00:54.39"><SPLITS/></RESULT><RESULT eventid="32" heatid="349" lane="3" points="150" resultid="2599" swimtime="00:01:47.02"><SPLITS><SPLIT distance="50" swimtime="00:00:50.90"/></SPLITS></RESULT><RESULT eventid="36" heatid="388" lane="3" points="150" resultid="2888" swimtime="00:00:41.85"><SPLITS/></RESULT><RESULT eventid="40" heatid="457" lane="3" points="153" resultid="3415" swimtime="00:01:27.46"><SPLITS><SPLIT distance="50" swimtime="00:00:41.42"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="233" birthdate="2014-01-01" firstname="Edoardo" gender="M" lastname="Dostetan Affuso" license="449618"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="31" lane="5" points="165" resultid="233" swimtime="00:00:47.30"><SPLITS/></RESULT><RESULT eventid="8" heatid="96" lane="3" points="200" resultid="720" swimtime="00:03:35.33"><SPLITS><SPLIT distance="50" swimtime="00:00:49.97"/><SPLIT distance="100" swimtime="00:01:44.49"/><SPLIT distance="150" swimtime="00:02:42.40"/></SPLITS></RESULT><RESULT eventid="10" heatid="140" lane="1" points="168" resultid="1052" swimtime="00:00:37.85"><SPLITS/></RESULT><RESULT eventid="12" heatid="176" lane="8" points="178" resultid="1335" swimtime="00:03:22.58"><SPLITS><SPLIT distance="50" swimtime="00:00:51.49"/><SPLIT distance="100" swimtime="00:01:43.41"/><SPLIT distance="150" swimtime="00:02:39.92"/></SPLITS></RESULT><RESULT eventid="26" heatid="251" lane="7" resultid="1861" swimtime="00:01:01.27"><SPLITS/></RESULT><RESULT eventid="30" heatid="313" lane="1" points="184" resultid="2327" swimtime="00:02:59.05"><SPLITS><SPLIT distance="50" swimtime="00:00:40.75"/><SPLIT distance="100" swimtime="00:01:26.59"/><SPLIT distance="150" swimtime="00:02:14.95"/></SPLITS></RESULT><RESULT eventid="32" heatid="348" lane="3" points="156" resultid="2592" swimtime="00:01:45.44"><SPLITS><SPLIT distance="50" swimtime="00:00:50.25"/></SPLITS></RESULT><RESULT eventid="40" heatid="459" lane="8" points="165" resultid="3436" swimtime="00:01:25.27"><SPLITS><SPLIT distance="50" swimtime="00:00:41.12"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="239" birthdate="2012-01-01" firstname="Bruno" gender="M" lastname="Matthes" license="445587"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="32" lane="3" points="156" resultid="239" swimtime="00:00:48.11"><SPLITS/></RESULT><RESULT eventid="8" heatid="96" lane="1" points="182" resultid="718" swimtime="00:03:42.23"><SPLITS><SPLIT distance="50" swimtime="00:00:48.86"/><SPLIT distance="100" swimtime="00:01:47.43"/><SPLIT distance="150" swimtime="00:02:47.72"/></SPLITS></RESULT><RESULT eventid="10" heatid="141" lane="3" points="190" resultid="1061" swimtime="00:00:36.34"><SPLITS/></RESULT><RESULT eventid="28" heatid="279" lane="2" points="154" resultid="2070" swimtime="00:00:44.15"><SPLITS/></RESULT><RESULT eventid="32" heatid="349" lane="7" points="153" resultid="2603" swimtime="00:01:46.13"><SPLITS><SPLIT distance="50" swimtime="00:00:49.34"/></SPLITS></RESULT><RESULT eventid="40" heatid="458" lane="4" points="192" resultid="3424" swimtime="00:01:21.16"><SPLITS><SPLIT distance="50" swimtime="00:00:37.67"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="247" birthdate="2012-01-01" firstname="Adrian" gender="M" lastname="Wyrwoll" license="421145"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="33" lane="3" points="130" resultid="247" swimtime="00:00:51.11"><SPLITS/></RESULT><RESULT eventid="6" heatid="75" lane="8" points="245" resultid="566" swimtime="00:01:18.93"><SPLITS><SPLIT distance="50" swimtime="00:00:36.93"/></SPLITS></RESULT><RESULT eventid="12" heatid="182" lane="8" points="253" resultid="1381" swimtime="00:03:00.04"><SPLITS><SPLIT distance="50" swimtime="00:00:36.94"/><SPLIT distance="100" swimtime="00:01:23.81"/><SPLIT distance="150" swimtime="00:02:19.14"/></SPLITS></RESULT><RESULT eventid="14" heatid="218" lane="3" points="206" resultid="1653" swimtime="00:01:27.25"><SPLITS><SPLIT distance="50" swimtime="00:00:42.32"/></SPLITS></RESULT><RESULT eventid="28" heatid="280" lane="1" points="209" resultid="2077" swimtime="00:00:39.94"><SPLITS/></RESULT><RESULT eventid="34" heatid="361" lane="2" points="243" resultid="2684" swimtime="00:02:56.80"><SPLITS><SPLIT distance="50" swimtime="00:00:39.55"/><SPLIT distance="100" swimtime="00:01:22.57"/><SPLIT distance="150" swimtime="00:02:11.03"/></SPLITS></RESULT><RESULT eventid="36" heatid="391" lane="5" points="239" resultid="2914" swimtime="00:00:35.84"><SPLITS/></RESULT><RESULT eventid="40" heatid="463" lane="6" points="254" resultid="3464" swimtime="00:01:13.99"><SPLITS><SPLIT distance="50" swimtime="00:00:35.52"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="265" birthdate="2011-01-01" firstname="Benedikt" gender="M" lastname="Deimling" license="483052"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="35" lane="7" points="204" resultid="265" swimtime="00:00:44.02"><SPLITS/></RESULT><RESULT eventid="8" heatid="98" lane="8" points="201" resultid="740" swimtime="00:03:34.74"><SPLITS><SPLIT distance="50" swimtime="00:00:46.22"/><SPLIT distance="100" swimtime="00:01:39.33"/><SPLIT distance="150" swimtime="00:02:38.42"/></SPLITS></RESULT><RESULT eventid="10" heatid="147" lane="1" points="256" resultid="1106" swimtime="00:00:32.93"><SPLITS/></RESULT><RESULT eventid="12" heatid="180" lane="4" points="240" resultid="1361" swimtime="00:03:03.21"><SPLITS><SPLIT distance="50" swimtime="00:00:38.10"/><SPLIT distance="100" swimtime="00:01:28.87"/><SPLIT distance="150" swimtime="00:02:22.59"/></SPLITS></RESULT><RESULT eventid="30" heatid="318" lane="3" points="278" resultid="2368" swimtime="00:02:36.10"><SPLITS><SPLIT distance="50" swimtime="00:00:35.51"/><SPLIT distance="100" swimtime="00:01:14.64"/><SPLIT distance="150" swimtime="00:01:56.06"/></SPLITS></RESULT><RESULT eventid="32" heatid="351" lane="6" points="188" resultid="2617" swimtime="00:01:39.13"><SPLITS><SPLIT distance="50" swimtime="00:00:45.84"/></SPLITS></RESULT><RESULT eventid="36" heatid="390" lane="8" points="204" resultid="2909" swimtime="00:00:37.81"><SPLITS/></RESULT><RESULT eventid="40" heatid="466" lane="8" points="303" resultid="3490" swimtime="00:01:09.76"><SPLITS><SPLIT distance="50" swimtime="00:00:33.95"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="272" birthdate="2012-01-01" firstname="Luis" gender="M" lastname="Alting van Geusau" license="435318"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="36" lane="6" points="307" resultid="272" swimtime="00:00:38.46"><SPLITS/></RESULT><RESULT eventid="8" heatid="99" lane="5" points="342" resultid="745" swimtime="00:03:00.01"><SPLITS><SPLIT distance="50" swimtime="00:00:43.27"/><SPLIT distance="100" swimtime="00:01:29.62"/><SPLIT distance="150" swimtime="00:02:16.59"/></SPLITS></RESULT><RESULT eventid="12" heatid="184" lane="1" points="345" resultid="1389" swimtime="00:02:42.47"><SPLITS><SPLIT distance="50" swimtime="00:00:36.51"/><SPLIT distance="100" swimtime="00:01:20.56"/><SPLIT distance="150" swimtime="00:02:05.24"/></SPLITS></RESULT><RESULT eventid="14" heatid="220" lane="4" points="272" resultid="1670" swimtime="00:01:19.57"><SPLITS><SPLIT distance="50" swimtime="00:00:38.42"/></SPLITS></RESULT><RESULT eventid="28" heatid="282" lane="7" points="293" resultid="2099" swimtime="00:00:35.67"><SPLITS/></RESULT><RESULT eventid="32" heatid="353" lane="1" points="315" resultid="2627" swimtime="00:01:23.53"><SPLITS><SPLIT distance="50" swimtime="00:00:40.25"/></SPLITS></RESULT><RESULT eventid="38" heatid="417" lane="6" points="294" resultid="3112" swimtime="00:02:48.25"><SPLITS><SPLIT distance="50" swimtime="00:00:38.96"/><SPLIT distance="100" swimtime="00:01:22.93"/><SPLIT distance="150" swimtime="00:02:04.94"/></SPLITS></RESULT><RESULT eventid="40" heatid="465" lane="6" points="347" resultid="3480" swimtime="00:01:06.63"><SPLITS><SPLIT distance="50" swimtime="00:00:32.00"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="286" birthdate="2010-01-01" firstname="Aurel" gender="M" lastname="Wyrwoll" license="421149"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="38" lane="4" points="425" resultid="286" swimtime="00:00:34.50"><SPLITS/></RESULT><RESULT eventid="8" heatid="93" lane="1" points="410" resultid="697" swimtime="00:02:49.46"><SPLITS><SPLIT distance="50" swimtime="00:00:36.90"/><SPLIT distance="100" swimtime="00:01:19.49"/><SPLIT distance="150" swimtime="00:02:05.59"/></SPLITS></RESULT><RESULT eventid="12" heatid="185" lane="7" points="327" resultid="1402" swimtime="00:02:45.42"><SPLITS><SPLIT distance="50" swimtime="00:00:39.18"/><SPLIT distance="100" swimtime="00:01:21.08"/><SPLIT distance="150" swimtime="00:02:05.06"/></SPLITS></RESULT><RESULT eventid="32" heatid="355" lane="8" points="423" resultid="2649" swimtime="00:01:15.73"><SPLITS><SPLIT distance="50" swimtime="00:00:35.30"/></SPLITS></RESULT><RESULT eventid="36" heatid="390" lane="3" points="267" resultid="2904" swimtime="00:00:34.55"><SPLITS/></RESULT><RESULT eventid="40" heatid="464" lane="4" points="314" resultid="3470" swimtime="00:01:08.89"><SPLITS><SPLIT distance="50" swimtime="00:00:31.68"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="305" birthdate="2009-01-01" firstname="Matteo" gender="M" lastname="Valtorta" license="392667"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="40" lane="7" resultid="305" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="4" heatid="62" lane="5" points="485" resultid="465" swimtime="00:04:40.03"><SPLITS><SPLIT distance="100" swimtime="00:01:06.60"/><SPLIT distance="200" swimtime="00:02:19.20"/><SPLIT distance="300" swimtime="00:03:32.03"/></SPLITS></RESULT><RESULT eventid="8" heatid="101" lane="8" points="421" resultid="763" swimtime="00:02:48.04"><SPLITS><SPLIT distance="50" swimtime="00:00:38.09"/><SPLIT distance="100" swimtime="00:01:20.33"/><SPLIT distance="150" swimtime="00:02:05.26"/></SPLITS></RESULT><RESULT eventid="10" heatid="153" lane="5" points="429" resultid="1158" swimtime="00:00:27.71"><SPLITS/></RESULT><RESULT eventid="18" heatid="233" lane="5" points="472" resultid="1756" swimtime="00:09:40.29"><SPLITS><SPLIT distance="100" swimtime="00:01:07.33"/><SPLIT distance="200" swimtime="00:02:20.48"/><SPLIT distance="300" swimtime="00:03:35.18"/><SPLIT distance="400" swimtime="00:04:50.38"/><SPLIT distance="500" swimtime="00:06:04.71"/><SPLIT distance="600" swimtime="00:07:17.85"/><SPLIT distance="700" swimtime="00:08:31.08"/></SPLITS></RESULT><RESULT eventid="30" heatid="325" lane="8" points="482" resultid="2425" swimtime="00:02:10.01"><SPLITS><SPLIT distance="50" swimtime="00:00:30.70"/><SPLIT distance="100" swimtime="00:01:03.87"/><SPLIT distance="150" swimtime="00:01:38.63"/></SPLITS></RESULT><RESULT eventid="32" heatid="356" lane="1" points="405" resultid="2650" swimtime="00:01:16.87"><SPLITS><SPLIT distance="50" swimtime="00:00:35.34"/></SPLITS></RESULT><RESULT eventid="40" heatid="471" lane="4" points="431" resultid="3525" swimtime="00:01:01.99"><SPLITS><SPLIT distance="50" swimtime="00:00:29.57"/></SPLITS></RESULT><RESULT eventid="42" heatid="481" lane="2" points="417" resultid="3592" swimtime="00:05:26.38"><SPLITS><SPLIT distance="50" swimtime="00:00:34.87"/><SPLIT distance="100" swimtime="00:01:15.44"/><SPLIT distance="150" swimtime="00:02:01.37"/><SPLIT distance="200" swimtime="00:02:43.68"/><SPLIT distance="250" swimtime="00:03:28.35"/><SPLIT distance="300" swimtime="00:04:14.04"/><SPLIT distance="350" swimtime="00:04:51.69"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="322" birthdate="2013-01-01" firstname="Magdalena" gender="F" lastname="Sirch" license="462118"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="43" lane="6" points="268" resultid="325" swimtime="00:06:06.52"><SPLITS><SPLIT distance="100" swimtime="00:01:26.61"/><SPLIT distance="200" swimtime="00:03:02.64"/><SPLIT distance="300" swimtime="00:04:36.71"/></SPLITS></RESULT><RESULT eventid="9" heatid="115" lane="1" points="284" resultid="865" swimtime="00:00:35.99"><SPLITS/></RESULT><RESULT eventid="11" heatid="160" lane="6" points="255" resultid="1208" swimtime="00:03:18.80"><SPLITS><SPLIT distance="50" swimtime="00:00:40.70"/><SPLIT distance="100" swimtime="00:01:31.73"/><SPLIT distance="150" swimtime="00:02:34.51"/></SPLITS></RESULT><RESULT eventid="23" heatid="241" lane="2" resultid="1793" swimtime="00:00:48.88"><SPLITS/></RESULT><RESULT eventid="29" heatid="296" lane="5" points="286" resultid="2202" swimtime="00:02:51.35"><SPLITS><SPLIT distance="50" swimtime="00:00:38.34"/><SPLIT distance="100" swimtime="00:01:22.19"/><SPLIT distance="150" swimtime="00:02:07.38"/></SPLITS></RESULT><RESULT eventid="31" heatid="334" lane="1" points="196" resultid="2483" swimtime="00:01:50.39"><SPLITS><SPLIT distance="50" swimtime="00:00:54.29"/></SPLITS></RESULT><RESULT eventid="35" heatid="367" lane="4" points="230" resultid="2730" swimtime="00:00:39.85"><SPLITS/></RESULT><RESULT eventid="39" heatid="431" lane="2" points="289" resultid="3211" swimtime="00:01:18.15"><SPLITS><SPLIT distance="50" swimtime="00:00:36.99"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="328" birthdate="2012-01-01" firstname="Antonia" gender="F" lastname="Lang" license="483067"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="44" lane="7" points="265" resultid="334" swimtime="00:06:08.03"><SPLITS><SPLIT distance="100" swimtime="00:01:24.65"/><SPLIT distance="200" swimtime="00:03:01.75"/><SPLIT distance="300" swimtime="00:04:37.72"/></SPLITS></RESULT><RESULT eventid="9" heatid="114" lane="7" points="307" resultid="863" swimtime="00:00:35.08"><SPLITS/></RESULT><RESULT eventid="13" heatid="199" lane="8" points="247" resultid="1511" swimtime="00:01:31.54"><SPLITS><SPLIT distance="50" swimtime="00:00:46.37"/></SPLITS></RESULT><RESULT eventid="27" heatid="262" lane="2" points="237" resultid="1941" swimtime="00:00:43.56"><SPLITS/></RESULT><RESULT eventid="29" heatid="295" lane="6" points="263" resultid="2195" swimtime="00:02:56.28"><SPLITS><SPLIT distance="50" swimtime="00:00:38.05"/><SPLIT distance="100" swimtime="00:01:24.28"/><SPLIT distance="150" swimtime="00:02:11.26"/></SPLITS></RESULT><RESULT eventid="37" heatid="405" lane="2" points="259" resultid="3016" swimtime="00:03:13.46"><SPLITS><SPLIT distance="50" swimtime="00:00:46.36"/><SPLIT distance="100" swimtime="00:01:36.75"/><SPLIT distance="150" swimtime="00:02:27.20"/></SPLITS></RESULT><RESULT comment="16:14 Start vor dem Startsignal" eventid="39" heatid="432" lane="5" resultid="3222" status="DSQ" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="332" birthdate="2012-01-01" firstname="Marlene" gender="F" lastname="Hambach" license="443546"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="45" lane="5" points="297" resultid="340" swimtime="00:05:54.27"><SPLITS><SPLIT distance="100" swimtime="00:01:23.38"/><SPLIT distance="200" swimtime="00:02:56.92"/><SPLIT distance="300" swimtime="00:04:30.02"/></SPLITS></RESULT><RESULT eventid="11" heatid="166" lane="6" points="305" resultid="1256" swimtime="00:03:07.30"><SPLITS><SPLIT distance="50" swimtime="00:00:43.41"/><SPLIT distance="100" swimtime="00:01:29.97"/><SPLIT distance="150" swimtime="00:02:25.66"/></SPLITS></RESULT><RESULT eventid="13" heatid="203" lane="8" points="349" resultid="1543" swimtime="00:01:21.57"><SPLITS><SPLIT distance="50" swimtime="00:00:40.19"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="340" birthdate="2013-01-01" firstname="Victoria" gender="F" lastname="Lucht" license="424870"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="47" lane="1" points="325" resultid="352" swimtime="00:05:43.53"><SPLITS><SPLIT distance="100" swimtime="00:01:23.21"/><SPLIT distance="200" swimtime="00:02:51.47"/><SPLIT distance="300" swimtime="00:04:20.16"/></SPLITS></RESULT><RESULT eventid="5" heatid="66" lane="1" points="312" resultid="489" swimtime="00:01:21.73"><SPLITS><SPLIT distance="50" swimtime="00:00:37.51"/></SPLITS></RESULT><RESULT eventid="11" heatid="169" lane="4" points="424" resultid="1278" swimtime="00:02:47.75"><SPLITS><SPLIT distance="50" swimtime="00:00:35.80"/><SPLIT distance="100" swimtime="00:01:17.85"/><SPLIT distance="150" swimtime="00:02:09.21"/></SPLITS></RESULT><RESULT eventid="13" heatid="204" lane="5" points="447" resultid="1548" swimtime="00:01:15.10"><SPLITS><SPLIT distance="50" swimtime="00:00:36.83"/></SPLITS></RESULT><RESULT eventid="19" heatid="235" lane="6" resultid="1767" swimtime="00:00:55.31"><SPLITS/></RESULT><RESULT eventid="27" heatid="268" lane="1" points="383" resultid="1988" swimtime="00:00:37.13"><SPLITS/></RESULT><RESULT eventid="33" heatid="358" lane="6" points="293" resultid="2665" swimtime="00:03:03.23"><SPLITS><SPLIT distance="50" swimtime="00:00:38.58"/><SPLIT distance="100" swimtime="00:01:24.58"/><SPLIT distance="150" swimtime="00:02:13.35"/></SPLITS></RESULT><RESULT eventid="37" heatid="409" lane="1" points="430" resultid="3047" swimtime="00:02:43.35"><SPLITS><SPLIT distance="50" swimtime="00:00:38.69"/><SPLIT distance="100" swimtime="00:01:20.23"/><SPLIT distance="150" swimtime="00:02:02.93"/></SPLITS></RESULT><RESULT eventid="39" heatid="437" lane="4" points="356" resultid="3261" swimtime="00:01:12.96"><SPLITS><SPLIT distance="50" swimtime="00:00:34.46"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="353" birthdate="2010-01-01" firstname="Louisa" gender="F" lastname="Seranski" license="419787"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="49" lane="4" points="368" resultid="370" swimtime="00:05:29.86"><SPLITS><SPLIT distance="100" swimtime="00:01:15.32"/><SPLIT distance="200" swimtime="00:02:39.47"/><SPLIT distance="300" swimtime="00:04:05.72"/></SPLITS></RESULT><RESULT eventid="9" heatid="122" lane="2" points="421" resultid="921" swimtime="00:00:31.56"><SPLITS/></RESULT><RESULT eventid="13" heatid="205" lane="8" points="396" resultid="1559" swimtime="00:01:18.23"><SPLITS><SPLIT distance="50" swimtime="00:00:39.13"/></SPLITS></RESULT><RESULT eventid="27" heatid="267" lane="4" points="399" resultid="1983" swimtime="00:00:36.63"><SPLITS/></RESULT><RESULT eventid="29" heatid="303" lane="7" points="388" resultid="2259" swimtime="00:02:34.82"><SPLITS><SPLIT distance="50" swimtime="00:00:35.72"/><SPLIT distance="100" swimtime="00:01:15.74"/><SPLIT distance="150" swimtime="00:01:55.92"/></SPLITS></RESULT><RESULT eventid="37" heatid="409" lane="3" points="419" resultid="3049" swimtime="00:02:44.81"><SPLITS><SPLIT distance="50" swimtime="00:00:39.59"/><SPLIT distance="100" swimtime="00:01:21.18"/><SPLIT distance="150" swimtime="00:02:03.47"/></SPLITS></RESULT><RESULT eventid="39" heatid="441" lane="8" points="392" resultid="3296" swimtime="00:01:10.62"><SPLITS><SPLIT distance="50" swimtime="00:00:34.43"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="361" birthdate="2009-01-01" firstname="Sandra" gender="F" lastname="Comteße" license="408110"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="50" lane="6" points="362" resultid="380" swimtime="00:05:31.59"><SPLITS><SPLIT distance="100" swimtime="00:01:15.23"/><SPLIT distance="200" swimtime="00:02:39.56"/><SPLIT distance="300" swimtime="00:04:05.87"/></SPLITS></RESULT><RESULT eventid="5" heatid="67" lane="2" points="317" resultid="498" swimtime="00:01:21.35"><SPLITS><SPLIT distance="50" swimtime="00:00:35.64"/></SPLITS></RESULT><RESULT eventid="11" heatid="168" lane="5" points="370" resultid="1271" swimtime="00:02:55.59"><SPLITS><SPLIT distance="50" swimtime="00:00:36.55"/><SPLIT distance="100" swimtime="00:01:21.50"/><SPLIT distance="150" swimtime="00:02:15.28"/></SPLITS></RESULT><RESULT eventid="15" heatid="226" lane="2" points="360" resultid="1713" swimtime="00:21:33.64"><SPLITS><SPLIT distance="100" swimtime="00:01:17.67"/><SPLIT distance="200" swimtime="00:02:42.49"/><SPLIT distance="300" swimtime="00:04:07.72"/><SPLIT distance="400" swimtime="00:05:32.34"/><SPLIT distance="500" swimtime="00:06:56.98"/><SPLIT distance="600" swimtime="00:08:22.54"/><SPLIT distance="700" swimtime="00:09:47.99"/><SPLIT distance="800" swimtime="00:11:14.11"/><SPLIT distance="900" swimtime="00:12:40.71"/><SPLIT distance="1000" swimtime="00:14:08.86"/><SPLIT distance="1100" swimtime="00:15:37.80"/><SPLIT distance="1200" swimtime="00:17:07.61"/><SPLIT distance="1300" swimtime="00:18:36.31"/><SPLIT distance="1400" swimtime="00:20:05.92"/></SPLITS></RESULT><RESULT eventid="29" heatid="303" lane="2" points="407" resultid="2254" swimtime="00:02:32.44"><SPLITS><SPLIT distance="50" swimtime="00:00:35.79"/><SPLIT distance="100" swimtime="00:01:14.35"/><SPLIT distance="150" swimtime="00:01:54.85"/></SPLITS></RESULT><RESULT eventid="35" heatid="376" lane="4" points="351" resultid="2801" swimtime="00:00:34.60"><SPLITS/></RESULT><RESULT eventid="37" heatid="408" lane="8" points="286" resultid="3046" swimtime="00:03:07.08"><SPLITS><SPLIT distance="50" swimtime="00:00:41.89"/><SPLIT distance="100" swimtime="00:01:26.59"/><SPLIT distance="150" swimtime="00:02:14.13"/></SPLITS></RESULT><RESULT eventid="39" heatid="444" lane="2" points="406" resultid="3314" swimtime="00:01:09.83"><SPLITS><SPLIT distance="50" swimtime="00:00:33.93"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="362" birthdate="2010-01-01" firstname="Lenya" gender="F" lastname="Horstmann" license="392670"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="50" lane="7" points="428" resultid="381" swimtime="00:05:13.59"><SPLITS><SPLIT distance="100" swimtime="00:01:12.42"/><SPLIT distance="200" swimtime="00:02:32.42"/></SPLITS></RESULT><RESULT eventid="5" heatid="68" lane="3" points="357" resultid="506" swimtime="00:01:18.15"><SPLITS><SPLIT distance="50" swimtime="00:00:36.06"/></SPLITS></RESULT><RESULT eventid="9" heatid="129" lane="7" points="522" resultid="981" swimtime="00:00:29.38"><SPLITS/></RESULT><RESULT eventid="11" heatid="170" lane="6" points="448" resultid="1288" swimtime="00:02:44.72"><SPLITS><SPLIT distance="50" swimtime="00:00:36.00"/><SPLIT distance="100" swimtime="00:01:19.17"/><SPLIT distance="150" swimtime="00:02:08.62"/></SPLITS></RESULT><RESULT eventid="27" heatid="270" lane="5" points="456" resultid="2007" swimtime="00:00:35.04"><SPLITS/></RESULT><RESULT eventid="29" heatid="303" lane="1" points="478" resultid="2253" swimtime="00:02:24.48"><SPLITS><SPLIT distance="50" swimtime="00:00:32.98"/><SPLIT distance="100" swimtime="00:01:08.98"/><SPLIT distance="150" swimtime="00:01:47.22"/></SPLITS></RESULT><RESULT eventid="35" heatid="379" lane="1" points="386" resultid="2820" swimtime="00:00:33.55"><SPLITS/></RESULT><RESULT eventid="39" heatid="448" lane="5" points="503" resultid="3347" swimtime="00:01:05.02"><SPLITS><SPLIT distance="50" swimtime="00:00:30.87"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="369" birthdate="2006-01-01" firstname="Ayla" gender="F" lastname="Hatil" license="348104"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="51" lane="7" points="457" resultid="388" swimtime="00:05:06.70"><SPLITS><SPLIT distance="100" swimtime="00:01:12.84"/><SPLIT distance="200" swimtime="00:02:30.37"/><SPLIT distance="300" swimtime="00:03:49.01"/></SPLITS></RESULT><RESULT eventid="7" heatid="92" lane="6" points="446" resultid="694" swimtime="00:03:01.82"><SPLITS><SPLIT distance="50" swimtime="00:00:41.89"/><SPLIT distance="100" swimtime="00:01:29.61"/><SPLIT distance="150" swimtime="00:02:15.76"/></SPLITS></RESULT><RESULT eventid="11" heatid="169" lane="6" points="434" resultid="1280" swimtime="00:02:46.57"><SPLITS><SPLIT distance="50" swimtime="00:00:35.48"/><SPLIT distance="100" swimtime="00:01:21.01"/><SPLIT distance="150" swimtime="00:02:07.69"/></SPLITS></RESULT><RESULT eventid="15" heatid="227" lane="2" points="475" resultid="1717" swimtime="00:19:39.59"><SPLITS><SPLIT distance="100" swimtime="00:01:16.46"/><SPLIT distance="200" swimtime="00:02:36.42"/><SPLIT distance="300" swimtime="00:03:56.30"/><SPLIT distance="400" swimtime="00:05:15.72"/><SPLIT distance="500" swimtime="00:06:35.02"/><SPLIT distance="600" swimtime="00:07:53.04"/><SPLIT distance="700" swimtime="00:09:11.68"/><SPLIT distance="800" swimtime="00:10:30.63"/><SPLIT distance="900" swimtime="00:11:49.56"/><SPLIT distance="1000" swimtime="00:13:08.51"/><SPLIT distance="1100" swimtime="00:14:26.63"/><SPLIT distance="1200" swimtime="00:15:45.00"/><SPLIT distance="1300" swimtime="00:17:03.65"/><SPLIT distance="1400" swimtime="00:18:22.06"/></SPLITS></RESULT><RESULT eventid="31" heatid="341" lane="4" points="429" resultid="2542" swimtime="00:01:24.97"><SPLITS><SPLIT distance="50" swimtime="00:00:39.94"/></SPLITS></RESULT><RESULT eventid="33" heatid="359" lane="7" points="306" resultid="2673" swimtime="00:03:00.57"><SPLITS><SPLIT distance="50" swimtime="00:00:39.78"/><SPLIT distance="100" swimtime="00:01:26.20"/><SPLIT distance="150" swimtime="00:02:15.25"/></SPLITS></RESULT><RESULT eventid="41" heatid="477" lane="6" points="453" resultid="3568" swimtime="00:05:46.69"><SPLITS><SPLIT distance="50" swimtime="00:00:36.17"/><SPLIT distance="100" swimtime="00:01:21.52"/><SPLIT distance="150" swimtime="00:02:08.07"/><SPLIT distance="200" swimtime="00:02:54.94"/><SPLIT distance="250" swimtime="00:03:41.76"/><SPLIT distance="300" swimtime="00:04:29.68"/><SPLIT distance="350" swimtime="00:05:08.76"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="377" birthdate="2007-01-01" firstname="Sophia" gender="F" lastname="Forster" license="363097"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="52" lane="7" points="497" resultid="396" swimtime="00:04:58.41"><SPLITS><SPLIT distance="100" swimtime="00:01:11.10"/><SPLIT distance="200" swimtime="00:02:27.41"/><SPLIT distance="300" swimtime="00:03:44.16"/></SPLITS></RESULT><RESULT eventid="7" heatid="92" lane="3" points="483" resultid="691" swimtime="00:02:57.04"><SPLITS><SPLIT distance="50" swimtime="00:00:41.20"/><SPLIT distance="100" swimtime="00:01:26.42"/><SPLIT distance="150" swimtime="00:02:12.56"/></SPLITS></RESULT><RESULT eventid="11" heatid="173" lane="2" points="456" resultid="1308" swimtime="00:02:43.78"><SPLITS><SPLIT distance="50" swimtime="00:00:35.64"/><SPLIT distance="100" swimtime="00:01:21.52"/><SPLIT distance="150" swimtime="00:02:07.39"/></SPLITS></RESULT><RESULT eventid="15" heatid="227" lane="6" points="478" resultid="1721" swimtime="00:19:36.84"><SPLITS><SPLIT distance="100" swimtime="00:01:16.30"/><SPLIT distance="200" swimtime="00:02:35.22"/><SPLIT distance="300" swimtime="00:03:54.30"/><SPLIT distance="400" swimtime="00:05:13.67"/><SPLIT distance="500" swimtime="00:06:33.53"/><SPLIT distance="600" swimtime="00:07:50.49"/><SPLIT distance="700" swimtime="00:09:08.90"/><SPLIT distance="800" swimtime="00:10:27.00"/><SPLIT distance="900" swimtime="00:11:46.17"/><SPLIT distance="1000" swimtime="00:13:05.71"/><SPLIT distance="1100" swimtime="00:14:24.30"/><SPLIT distance="1200" swimtime="00:15:42.94"/><SPLIT distance="1300" swimtime="00:17:01.80"/><SPLIT distance="1400" swimtime="00:18:20.11"/></SPLITS></RESULT><RESULT eventid="31" heatid="342" lane="8" points="384" resultid="2554" swimtime="00:01:28.17"><SPLITS><SPLIT distance="50" swimtime="00:00:42.59"/></SPLITS></RESULT><RESULT eventid="33" heatid="359" lane="3" points="380" resultid="2669" swimtime="00:02:48.05"><SPLITS><SPLIT distance="50" swimtime="00:00:37.92"/><SPLIT distance="100" swimtime="00:01:18.94"/><SPLIT distance="150" swimtime="00:02:02.58"/></SPLITS></RESULT><RESULT eventid="41" heatid="478" lane="5" points="500" resultid="3574" swimtime="00:05:35.38"><SPLITS><SPLIT distance="50" swimtime="00:00:35.34"/><SPLIT distance="100" swimtime="00:01:16.38"/><SPLIT distance="200" swimtime="00:02:47.39"/><SPLIT distance="250" swimtime="00:03:33.43"/><SPLIT distance="300" swimtime="00:04:19.06"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="379" birthdate="2013-01-01" firstname="Edoardo" gender="M" lastname="Lepore" license="483064"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="53" lane="3" points="111" resultid="399" swimtime="00:07:37.54"><SPLITS><SPLIT distance="100" swimtime="00:01:45.22"/><SPLIT distance="200" swimtime="00:03:43.47"/><SPLIT distance="300" swimtime="00:05:45.07"/></SPLITS></RESULT><RESULT eventid="10" heatid="138" lane="1" points="133" resultid="1037" swimtime="00:00:40.89"><SPLITS/></RESULT><RESULT eventid="12" heatid="175" lane="6" points="137" resultid="1327" swimtime="00:03:40.97"><SPLITS><SPLIT distance="50" swimtime="00:02:50.39"/><SPLIT distance="100" swimtime="00:01:46.62"/><SPLIT distance="150" swimtime="00:02:50.39"/></SPLITS></RESULT><RESULT eventid="14" heatid="212" lane="3" points="125" resultid="1607" swimtime="00:01:43.03"><SPLITS><SPLIT distance="50" swimtime="00:00:51.21"/></SPLITS></RESULT><RESULT eventid="20" heatid="236" lane="7" resultid="1775" swimtime="00:01:12.60"><SPLITS/></RESULT><RESULT eventid="24" heatid="244" lane="3" resultid="1816" swimtime="00:01:01.14"><SPLITS/></RESULT><RESULT eventid="30" heatid="311" lane="1" points="109" resultid="2312" swimtime="00:03:33.31"><SPLITS><SPLIT distance="50" swimtime="00:00:48.12"/><SPLIT distance="100" swimtime="00:01:43.59"/><SPLIT distance="150" swimtime="00:02:41.26"/></SPLITS></RESULT><RESULT comment="14:25 Der Sportler führte mehrere Wechselbeinschläge aus" eventid="36" heatid="384" lane="8" resultid="2862" status="DSQ" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="40" heatid="455" lane="7" points="108" resultid="3404" swimtime="00:01:38.20"><SPLITS><SPLIT distance="50" swimtime="00:00:45.51"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="385" birthdate="2015-01-01" firstname="Moritz" gender="M" lastname="Fink" license="489624"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="54" lane="6" points="184" resultid="407" swimtime="00:06:26.59"><SPLITS><SPLIT distance="100" swimtime="00:01:24.94"/><SPLIT distance="200" swimtime="00:03:05.37"/><SPLIT distance="300" swimtime="00:04:47.16"/></SPLITS></RESULT><RESULT eventid="10" heatid="140" lane="6" points="194" resultid="1057" swimtime="00:00:36.11"><SPLITS/></RESULT><RESULT eventid="12" heatid="175" lane="5" points="140" resultid="1326" swimtime="00:03:39.49"><SPLITS><SPLIT distance="50" swimtime="00:00:53.05"/><SPLIT distance="100" swimtime="00:01:47.51"/><SPLIT distance="150" swimtime="00:02:55.30"/></SPLITS></RESULT><RESULT eventid="14" heatid="212" lane="4" points="126" resultid="1608" swimtime="00:01:42.69"><SPLITS><SPLIT distance="50" swimtime="00:00:48.28"/></SPLITS></RESULT><RESULT eventid="30" heatid="312" lane="4" points="187" resultid="2322" swimtime="00:02:58.33"><SPLITS><SPLIT distance="50" swimtime="00:00:38.26"/><SPLIT distance="100" swimtime="00:01:25.24"/><SPLIT distance="150" swimtime="00:02:13.44"/></SPLITS></RESULT><RESULT eventid="36" heatid="385" lane="7" points="87" resultid="2869" swimtime="00:00:50.23"><SPLITS/></RESULT><RESULT comment="15:36 Der Sportler hat nach dem erlaubten Armzug in Bauchlage die 100m Wende nicht unverzüglich eingeleitet" eventid="38" heatid="414" lane="8" resultid="3090" status="DSQ" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="40" heatid="457" lane="5" points="181" resultid="3417" swimtime="00:01:22.72"><SPLITS><SPLIT distance="50" swimtime="00:00:38.96"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="397" birthdate="2013-01-01" firstname="Miron" gender="M" lastname="Voinov" license="446393"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="56" lane="6" points="211" resultid="423" swimtime="00:06:09.47"><SPLITS><SPLIT distance="100" swimtime="00:01:22.54"/><SPLIT distance="200" swimtime="00:02:59.75"/><SPLIT distance="300" swimtime="00:04:37.66"/></SPLITS></RESULT><RESULT eventid="10" heatid="143" lane="6" points="217" resultid="1079" swimtime="00:00:34.77"><SPLITS/></RESULT><RESULT eventid="12" heatid="177" lane="5" points="166" resultid="1339" swimtime="00:03:27.28"><SPLITS><SPLIT distance="50" swimtime="00:00:49.91"/><SPLIT distance="100" swimtime="00:01:39.45"/><SPLIT distance="150" swimtime="00:02:42.91"/></SPLITS></RESULT><RESULT eventid="14" heatid="220" lane="3" points="224" resultid="1669" swimtime="00:01:24.94"><SPLITS><SPLIT distance="50" swimtime="00:00:41.74"/></SPLITS></RESULT><RESULT eventid="20" heatid="236" lane="3" resultid="1771" swimtime="00:00:49.20"><SPLITS/></RESULT><RESULT eventid="24" heatid="245" lane="6" resultid="1825" swimtime="00:00:46.26"><SPLITS/></RESULT><RESULT eventid="32" heatid="349" lane="1" points="156" resultid="2597" swimtime="00:01:45.66"><SPLITS><SPLIT distance="50" swimtime="00:00:51.28"/></SPLITS></RESULT><RESULT eventid="38" heatid="416" lane="4" points="228" resultid="3102" swimtime="00:03:02.96"><SPLITS><SPLIT distance="50" swimtime="00:00:42.90"/><SPLIT distance="100" swimtime="00:01:29.56"/><SPLIT distance="150" swimtime="00:02:17.68"/></SPLITS></RESULT><RESULT eventid="40" heatid="462" lane="5" points="234" resultid="3456" swimtime="00:01:16.04"><SPLITS><SPLIT distance="50" swimtime="00:00:35.96"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="422" birthdate="2010-01-01" firstname="Lennart Matthias" gender="M" lastname="Schlobach" license="462467"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="60" lane="3" points="454" resultid="451" swimtime="00:04:46.22"><SPLITS><SPLIT distance="100" swimtime="00:01:08.15"/><SPLIT distance="200" swimtime="00:02:21.00"/><SPLIT distance="300" swimtime="00:03:34.22"/></SPLITS></RESULT><RESULT eventid="6" heatid="76" lane="2" points="373" resultid="568" swimtime="00:01:08.69"><SPLITS><SPLIT distance="50" swimtime="00:00:32.47"/></SPLITS></RESULT><RESULT eventid="12" heatid="186" lane="1" points="411" resultid="1404" swimtime="00:02:33.27"><SPLITS><SPLIT distance="50" swimtime="00:00:33.05"/><SPLIT distance="100" swimtime="00:01:13.14"/><SPLIT distance="150" swimtime="00:02:00.11"/></SPLITS></RESULT><RESULT eventid="14" heatid="222" lane="5" points="367" resultid="1686" swimtime="00:01:12.03"><SPLITS><SPLIT distance="50" swimtime="00:00:35.90"/></SPLITS></RESULT><RESULT eventid="18" heatid="233" lane="2" points="450" resultid="1754" swimtime="00:09:49.68"><SPLITS><SPLIT distance="100" swimtime="00:01:10.14"/><SPLIT distance="200" swimtime="00:02:24.16"/><SPLIT distance="300" swimtime="00:03:38.16"/><SPLIT distance="400" swimtime="00:04:52.36"/><SPLIT distance="500" swimtime="00:06:06.98"/><SPLIT distance="600" swimtime="00:07:21.47"/><SPLIT distance="700" swimtime="00:08:36.42"/></SPLITS></RESULT><RESULT eventid="30" heatid="322" lane="3" points="461" resultid="2398" swimtime="00:02:12.02"><SPLITS><SPLIT distance="50" swimtime="00:00:30.74"/><SPLIT distance="100" swimtime="00:01:04.06"/><SPLIT distance="150" swimtime="00:01:38.91"/></SPLITS></RESULT><RESULT eventid="34" heatid="361" lane="4" points="346" resultid="2685" swimtime="00:02:37.11"><SPLITS><SPLIT distance="50" swimtime="00:00:34.83"/><SPLIT distance="100" swimtime="00:01:16.40"/><SPLIT distance="150" swimtime="00:01:57.51"/></SPLITS></RESULT><RESULT eventid="38" heatid="418" lane="3" points="377" resultid="3116" swimtime="00:02:34.89"><SPLITS><SPLIT distance="50" swimtime="00:00:37.72"/><SPLIT distance="100" swimtime="00:01:16.50"/><SPLIT distance="150" swimtime="00:01:56.52"/></SPLITS></RESULT><RESULT eventid="42" heatid="480" lane="3" points="439" resultid="3587" swimtime="00:05:20.64"><SPLITS><SPLIT distance="50" swimtime="00:00:33.94"/><SPLIT distance="100" swimtime="00:01:14.65"/><SPLIT distance="150" swimtime="00:01:55.65"/><SPLIT distance="200" swimtime="00:02:35.35"/><SPLIT distance="250" swimtime="00:03:24.03"/><SPLIT distance="300" swimtime="00:04:12.29"/><SPLIT distance="350" swimtime="00:04:46.83"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="431" birthdate="2011-01-01" firstname="Edouard" gender="M" lastname="Plantet-Vuc" license="453053"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="61" lane="6" points="443" resultid="460" swimtime="00:04:48.50"><SPLITS><SPLIT distance="100" swimtime="00:01:11.58"/><SPLIT distance="200" swimtime="00:02:25.51"/><SPLIT distance="300" swimtime="00:03:37.78"/></SPLITS></RESULT><RESULT eventid="8" heatid="100" lane="1" points="354" resultid="749" swimtime="00:02:58.02"><SPLITS><SPLIT distance="50" swimtime="00:00:40.41"/><SPLIT distance="100" swimtime="00:01:26.95"/><SPLIT distance="150" swimtime="00:02:11.90"/></SPLITS></RESULT><RESULT eventid="12" heatid="187" lane="1" points="363" resultid="1412" swimtime="00:02:39.78"><SPLITS><SPLIT distance="50" swimtime="00:00:37.16"/><SPLIT distance="100" swimtime="00:01:18.11"/><SPLIT distance="150" swimtime="00:02:04.57"/></SPLITS></RESULT><RESULT eventid="14" heatid="222" lane="4" points="321" resultid="1685" swimtime="00:01:15.36"><SPLITS><SPLIT distance="50" swimtime="00:00:36.59"/></SPLITS></RESULT><RESULT eventid="18" heatid="232" lane="4" points="440" resultid="1750" swimtime="00:09:54.28"><SPLITS><SPLIT distance="100" swimtime="00:01:12.31"/><SPLIT distance="200" swimtime="00:02:28.20"/><SPLIT distance="300" swimtime="00:03:44.31"/><SPLIT distance="400" swimtime="00:04:58.90"/><SPLIT distance="500" swimtime="00:06:13.76"/><SPLIT distance="600" swimtime="00:07:28.35"/><SPLIT distance="700" swimtime="00:08:41.73"/></SPLITS></RESULT><RESULT eventid="30" heatid="322" lane="5" points="435" resultid="2400" swimtime="00:02:14.61"><SPLITS><SPLIT distance="50" swimtime="00:00:32.09"/><SPLIT distance="100" swimtime="00:01:05.67"/><SPLIT distance="150" swimtime="00:01:40.69"/></SPLITS></RESULT><RESULT eventid="32" heatid="352" lane="6" points="305" resultid="2624" swimtime="00:01:24.49"><SPLITS><SPLIT distance="50" swimtime="00:00:40.13"/></SPLITS></RESULT><RESULT eventid="38" heatid="418" lane="6" points="365" resultid="3118" swimtime="00:02:36.54"><SPLITS><SPLIT distance="50" swimtime="00:00:37.36"/><SPLIT distance="100" swimtime="00:01:17.51"/><SPLIT distance="150" swimtime="00:01:57.34"/></SPLITS></RESULT><RESULT eventid="42" heatid="480" lane="7" points="388" resultid="3590" swimtime="00:05:34.27"><SPLITS><SPLIT distance="50" swimtime="00:00:36.45"/><SPLIT distance="100" swimtime="00:01:22.02"/><SPLIT distance="150" swimtime="00:02:04.48"/><SPLIT distance="200" swimtime="00:02:45.95"/><SPLIT distance="250" swimtime="00:03:33.19"/><SPLIT distance="300" swimtime="00:04:21.08"/><SPLIT distance="350" swimtime="00:04:58.08"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="454" birthdate="2008-01-01" firstname="Lilly" gender="F" lastname="Zöckler" license="414291"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="5" heatid="68" lane="2" points="383" resultid="505" swimtime="00:01:16.33"><SPLITS><SPLIT distance="50" swimtime="00:00:35.46"/></SPLITS></RESULT><RESULT eventid="9" heatid="127" lane="6" points="409" resultid="964" swimtime="00:00:31.88"><SPLITS/></RESULT><RESULT eventid="11" heatid="170" lane="2" points="392" resultid="1284" swimtime="00:02:52.24"><SPLITS><SPLIT distance="50" swimtime="00:00:34.87"/><SPLIT distance="100" swimtime="00:01:24.09"/><SPLIT distance="150" swimtime="00:02:12.95"/></SPLITS></RESULT><RESULT eventid="29" heatid="304" lane="1" points="407" resultid="2261" swimtime="00:02:32.34"><SPLITS><SPLIT distance="50" swimtime="00:00:34.96"/><SPLIT distance="100" swimtime="00:01:13.49"/><SPLIT distance="150" swimtime="00:01:54.55"/></SPLITS></RESULT><RESULT eventid="31" heatid="341" lane="2" points="391" resultid="2540" swimtime="00:01:27.67"><SPLITS><SPLIT distance="50" swimtime="00:00:41.85"/></SPLITS></RESULT><RESULT eventid="35" heatid="376" lane="5" points="390" resultid="2802" swimtime="00:00:33.43"><SPLITS/></RESULT><RESULT eventid="39" heatid="447" lane="7" points="417" resultid="3341" swimtime="00:01:09.17"><SPLITS><SPLIT distance="50" swimtime="00:00:32.82"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="455" birthdate="2007-01-01" firstname="Anna" gender="F" lastname="Dinkel" license="367689"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="5" heatid="68" lane="5" points="404" resultid="508" swimtime="00:01:15.03"><SPLITS><SPLIT distance="50" swimtime="00:00:34.69"/></SPLITS></RESULT><RESULT eventid="11" heatid="174" lane="1" points="470" resultid="1315" swimtime="00:02:42.12"><SPLITS><SPLIT distance="50" swimtime="00:00:37.14"/><SPLIT distance="100" swimtime="00:01:16.96"/><SPLIT distance="150" swimtime="00:02:04.77"/></SPLITS></RESULT><RESULT eventid="13" heatid="208" lane="3" points="427" resultid="1577" swimtime="00:01:16.26"><SPLITS><SPLIT distance="50" swimtime="00:00:37.15"/></SPLITS></RESULT><RESULT eventid="27" heatid="271" lane="8" points="405" resultid="2017" swimtime="00:00:36.45"><SPLITS/></RESULT><RESULT eventid="33" heatid="360" lane="1" points="389" resultid="2675" swimtime="00:02:46.84"><SPLITS><SPLIT distance="50" swimtime="00:00:37.22"/><SPLIT distance="100" swimtime="00:01:18.48"/><SPLIT distance="150" swimtime="00:02:04.00"/></SPLITS></RESULT><RESULT eventid="37" heatid="411" lane="4" points="452" resultid="3066" swimtime="00:02:40.72"><SPLITS><SPLIT distance="100" swimtime="00:01:17.79"/></SPLITS></RESULT><RESULT eventid="41" heatid="478" lane="7" points="445" resultid="3576" swimtime="00:05:48.78"><SPLITS><SPLIT distance="50" swimtime="00:00:36.78"/><SPLIT distance="100" swimtime="00:01:22.85"/><SPLIT distance="150" swimtime="00:02:07.57"/><SPLIT distance="200" swimtime="00:02:50.83"/><SPLIT distance="250" swimtime="00:03:39.24"/><SPLIT distance="300" swimtime="00:04:28.64"/><SPLIT distance="350" swimtime="00:05:09.21"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="459" birthdate="2006-01-01" firstname="Sophia" gender="F" lastname="Horstmann" license="344033"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="5" heatid="70" lane="3" points="472" resultid="522" swimtime="00:01:11.25"><SPLITS><SPLIT distance="50" swimtime="00:00:33.65"/></SPLITS></RESULT><RESULT eventid="11" heatid="171" lane="1" points="519" resultid="1291" swimtime="00:02:36.93"><SPLITS><SPLIT distance="50" swimtime="00:00:33.52"/><SPLIT distance="100" swimtime="00:01:15.91"/><SPLIT distance="150" swimtime="00:02:03.32"/></SPLITS></RESULT><RESULT eventid="13" heatid="209" lane="1" points="505" resultid="1583" swimtime="00:01:12.14"><SPLITS><SPLIT distance="50" swimtime="00:00:35.74"/></SPLITS></RESULT><RESULT eventid="27" heatid="272" lane="5" points="543" resultid="2022" swimtime="00:00:33.07"><SPLITS/></RESULT><RESULT eventid="29" heatid="305" lane="5" points="558" resultid="2271" swimtime="00:02:17.21"><SPLITS><SPLIT distance="50" swimtime="00:00:31.95"/><SPLIT distance="100" swimtime="00:01:07.54"/><SPLIT distance="150" swimtime="00:01:43.63"/></SPLITS></RESULT><RESULT eventid="35" heatid="382" lane="7" points="504" resultid="2850" swimtime="00:00:30.68"><SPLITS/></RESULT><RESULT eventid="37" heatid="412" lane="3" points="517" resultid="3073" swimtime="00:02:33.66"><SPLITS><SPLIT distance="100" swimtime="00:01:15.53"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="467" birthdate="2008-01-01" firstname="Elena" gender="F" lastname="Harteneck" license="392664"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="5" heatid="71" lane="7" points="480" resultid="534" swimtime="00:01:10.85"><SPLITS><SPLIT distance="50" swimtime="00:00:31.69"/></SPLITS></RESULT><RESULT eventid="9" heatid="129" lane="3" points="510" resultid="977" swimtime="00:00:29.61"><SPLITS/></RESULT><RESULT eventid="13" heatid="206" lane="4" points="430" resultid="1563" swimtime="00:01:16.11"><SPLITS><SPLIT distance="50" swimtime="00:00:37.00"/></SPLITS></RESULT><RESULT eventid="29" heatid="304" lane="3" points="492" resultid="2263" swimtime="00:02:23.04"><SPLITS><SPLIT distance="50" swimtime="00:00:33.45"/><SPLIT distance="100" swimtime="00:01:09.61"/><SPLIT distance="150" swimtime="00:01:47.77"/></SPLITS></RESULT><RESULT eventid="33" heatid="360" lane="7" points="400" resultid="2681" swimtime="00:02:45.21"><SPLITS><SPLIT distance="50" swimtime="00:00:35.10"/><SPLIT distance="100" swimtime="00:01:16.82"/><SPLIT distance="150" swimtime="00:02:00.58"/></SPLITS></RESULT><RESULT eventid="35" heatid="380" lane="4" points="435" resultid="2831" swimtime="00:00:32.22"><SPLITS/></RESULT><RESULT eventid="39" heatid="450" lane="3" points="558" resultid="3360" swimtime="00:01:02.78"><SPLITS><SPLIT distance="50" swimtime="00:00:30.34"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="491" birthdate="2007-01-01" firstname="Gregor" gender="M" lastname="Comteße" license="409328"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="6" heatid="77" lane="5" points="386" resultid="579" swimtime="00:01:07.87"><SPLITS><SPLIT distance="50" swimtime="00:00:30.50"/></SPLITS></RESULT><RESULT eventid="10" heatid="152" lane="5" points="472" resultid="1150" swimtime="00:00:26.84"><SPLITS/></RESULT><RESULT eventid="12" heatid="188" lane="6" points="445" resultid="1425" swimtime="00:02:29.28"><SPLITS><SPLIT distance="50" swimtime="00:00:31.15"/><SPLIT distance="100" swimtime="00:01:10.74"/><SPLIT distance="150" swimtime="00:01:56.65"/></SPLITS></RESULT><RESULT eventid="30" heatid="325" lane="6" points="493" resultid="2423" swimtime="00:02:09.07"><SPLITS><SPLIT distance="50" swimtime="00:00:29.71"/><SPLIT distance="100" swimtime="00:01:02.79"/><SPLIT distance="150" swimtime="00:01:36.65"/></SPLITS></RESULT><RESULT eventid="40" heatid="475" lane="7" points="427" resultid="3558" swimtime="00:01:02.21"><SPLITS><SPLIT distance="50" swimtime="00:00:28.75"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="508" birthdate="2009-01-01" firstname="Mathilda" gender="F" lastname="Wery" license="381312"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="7" heatid="91" lane="3" points="492" resultid="683" swimtime="00:02:55.98"><SPLITS><SPLIT distance="50" swimtime="00:00:39.45"/><SPLIT distance="100" swimtime="00:01:24.51"/><SPLIT distance="150" swimtime="00:02:10.48"/></SPLITS></RESULT><RESULT eventid="11" heatid="174" lane="3" points="543" resultid="1317" swimtime="00:02:34.53"><SPLITS><SPLIT distance="50" swimtime="00:00:33.60"/><SPLIT distance="100" swimtime="00:01:11.99"/><SPLIT distance="150" swimtime="00:01:58.18"/></SPLITS></RESULT><RESULT eventid="13" heatid="209" lane="2" points="515" resultid="1584" swimtime="00:01:11.65"><SPLITS><SPLIT distance="50" swimtime="00:00:35.11"/></SPLITS></RESULT><RESULT eventid="27" heatid="272" lane="7" points="523" resultid="2023" swimtime="00:00:33.48"><SPLITS/></RESULT><RESULT eventid="31" heatid="343" lane="4" points="486" resultid="2558" swimtime="00:01:21.55"><SPLITS><SPLIT distance="50" swimtime="00:00:37.92"/></SPLITS></RESULT><RESULT eventid="37" heatid="412" lane="4" points="536" resultid="3074" swimtime="00:02:31.82"><SPLITS><SPLIT distance="100" swimtime="00:01:13.97"/></SPLITS></RESULT><RESULT eventid="41" heatid="478" lane="2" points="528" resultid="3571" swimtime="00:05:29.35"><SPLITS><SPLIT distance="50" swimtime="00:00:34.16"/><SPLIT distance="100" swimtime="00:01:15.45"/><SPLIT distance="150" swimtime="00:01:56.96"/><SPLIT distance="200" swimtime="00:02:38.30"/><SPLIT distance="250" swimtime="00:03:25.55"/><SPLIT distance="300" swimtime="00:04:13.90"/><SPLIT distance="350" swimtime="00:04:52.01"/></SPLITS></RESULT></RESULTS></ATHLETE></ATHLETES><RELAYS/></CLUB><CLUB code="4529" name="TV Münchberg" nation="GER" region="02" shortname="Münchber" type="CLUB"><CONTACT city="Münchberg" country="GER" email="nicole.hertrich94@gmail.com" name="Wagner, Nicole" phone="09251/8507780" street="Bayreuther Str. 62" zip="95213"/><OFFICIALS/><ATHLETES><ATHLETE athleteid="33" birthdate="2016-01-01" firstname="Marie" gender="F" lastname="Dillner" license="485588"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="5" lane="5" points="141" resultid="33" swimtime="00:00:56.19"><SPLITS/></RESULT><RESULT eventid="9" heatid="108" lane="6" points="164" resultid="814" swimtime="00:00:43.17"><SPLITS/></RESULT><RESULT eventid="29" heatid="288" lane="5" points="155" resultid="2141" swimtime="00:03:30.27"><SPLITS><SPLIT distance="50" swimtime="00:00:44.17"/><SPLIT distance="100" swimtime="00:01:40.39"/><SPLIT distance="150" swimtime="00:02:37.07"/></SPLITS></RESULT><RESULT eventid="31" heatid="329" lane="1" points="132" resultid="2443" swimtime="00:02:05.69"><SPLITS><SPLIT distance="50" swimtime="00:01:00.45"/></SPLITS></RESULT><RESULT eventid="39" heatid="424" lane="3" points="141" resultid="3157" swimtime="00:01:39.13"><SPLITS><SPLIT distance="50" swimtime="00:00:46.18"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="193" birthdate="2016-01-01" firstname="Benedikt" gender="M" lastname="Ramming" license="485592"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="26" lane="4" points="80" resultid="193" swimtime="00:01:00.02"><SPLITS/></RESULT><RESULT eventid="10" heatid="135" lane="3" points="97" resultid="1015" swimtime="00:00:45.37"><SPLITS/></RESULT><RESULT eventid="14" heatid="210" lane="6" points="85" resultid="1595" swimtime="00:01:56.98"><SPLITS><SPLIT distance="50" swimtime="00:00:57.11"/></SPLITS></RESULT><RESULT eventid="28" heatid="275" lane="1" points="84" resultid="2039" swimtime="00:00:54.13"><SPLITS/></RESULT><RESULT eventid="30" heatid="309" lane="5" points="85" resultid="2300" swimtime="00:03:51.70"><SPLITS><SPLIT distance="50" swimtime="00:00:53.32"/><SPLIT distance="100" swimtime="00:01:56.38"/><SPLIT distance="150" swimtime="00:02:55.16"/></SPLITS></RESULT><RESULT eventid="36" heatid="383" lane="3" points="58" resultid="2852" swimtime="00:00:57.48"><SPLITS/></RESULT><RESULT eventid="40" heatid="453" lane="4" points="99" resultid="3385" swimtime="00:01:40.97"><SPLITS><SPLIT distance="50" swimtime="00:00:49.13"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="313" birthdate="2014-01-01" firstname="Emma" gender="F" lastname="Skaper" license="462940"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="42" lane="3" points="295" resultid="314" swimtime="00:05:54.78"><SPLITS><SPLIT distance="100" swimtime="00:01:21.84"/><SPLIT distance="200" swimtime="00:02:54.31"/><SPLIT distance="300" swimtime="00:04:27.23"/></SPLITS></RESULT><RESULT eventid="7" heatid="83" lane="6" points="283" resultid="623" swimtime="00:03:31.46"><SPLITS><SPLIT distance="50" swimtime="00:00:48.94"/><SPLIT distance="100" swimtime="00:01:44.14"/><SPLIT distance="150" swimtime="00:02:38.45"/></SPLITS></RESULT><RESULT eventid="11" heatid="163" lane="2" points="286" resultid="1228" swimtime="00:03:11.21"><SPLITS><SPLIT distance="50" swimtime="00:00:44.51"/><SPLIT distance="100" swimtime="00:01:33.28"/><SPLIT distance="150" swimtime="00:02:30.58"/></SPLITS></RESULT><RESULT eventid="13" heatid="198" lane="5" points="235" resultid="1500" swimtime="00:01:33.01"><SPLITS/></RESULT><RESULT eventid="29" heatid="296" lane="7" points="315" resultid="2204" swimtime="00:02:45.92"><SPLITS><SPLIT distance="50" swimtime="00:00:36.97"/><SPLIT distance="100" swimtime="00:01:19.99"/><SPLIT distance="150" swimtime="00:02:03.45"/></SPLITS></RESULT><RESULT eventid="33" heatid="358" lane="7" points="194" resultid="2666" swimtime="00:03:30.34"><SPLITS><SPLIT distance="50" swimtime="00:00:45.64"/><SPLIT distance="100" swimtime="00:01:39.79"/><SPLIT distance="150" swimtime="00:02:37.04"/></SPLITS></RESULT><RESULT eventid="39" heatid="432" lane="2" points="290" resultid="3219" swimtime="00:01:18.11"><SPLITS><SPLIT distance="50" swimtime="00:00:37.88"/></SPLITS></RESULT><RESULT eventid="41" heatid="476" lane="5" points="293" resultid="3562" swimtime="00:06:40.61"><SPLITS><SPLIT distance="50" swimtime="00:00:45.19"/><SPLIT distance="100" swimtime="00:01:38.21"/><SPLIT distance="150" swimtime="00:02:30.10"/><SPLIT distance="200" swimtime="00:03:20.35"/><SPLIT distance="250" swimtime="00:04:14.99"/><SPLIT distance="300" swimtime="00:05:10.91"/><SPLIT distance="350" swimtime="00:05:57.59"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="447" birthdate="2013-01-01" firstname="Theresa" gender="F" lastname="Fischer" license="463322"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="5" heatid="65" lane="7" points="210" resultid="487" swimtime="00:01:33.28"><SPLITS><SPLIT distance="50" swimtime="00:00:40.94"/></SPLITS></RESULT><RESULT eventid="11" heatid="162" lane="4" points="249" resultid="1222" swimtime="00:03:20.45"><SPLITS><SPLIT distance="50" swimtime="00:00:42.80"/><SPLIT distance="100" swimtime="00:01:35.13"/><SPLIT distance="150" swimtime="00:02:35.67"/></SPLITS></RESULT><RESULT eventid="13" heatid="197" lane="2" points="227" resultid="1489" swimtime="00:01:34.17"><SPLITS><SPLIT distance="50" swimtime="00:00:46.17"/></SPLITS></RESULT><RESULT eventid="33" heatid="358" lane="1" points="200" resultid="2661" swimtime="00:03:28.29"><SPLITS><SPLIT distance="50" swimtime="00:00:46.72"/><SPLIT distance="100" swimtime="00:01:39.96"/><SPLIT distance="150" swimtime="00:02:38.00"/></SPLITS></RESULT><RESULT eventid="35" heatid="372" lane="3" points="240" resultid="2769" swimtime="00:00:39.28"><SPLITS/></RESULT><RESULT eventid="41" heatid="476" lane="3" points="258" resultid="3560" swimtime="00:06:58.05"><SPLITS><SPLIT distance="50" swimtime="00:00:46.52"/><SPLIT distance="100" swimtime="00:01:41.36"/><SPLIT distance="150" swimtime="00:02:35.67"/><SPLIT distance="200" swimtime="00:03:28.98"/><SPLIT distance="250" swimtime="00:04:28.19"/><SPLIT distance="300" swimtime="00:05:30.14"/><SPLIT distance="350" swimtime="00:06:17.92"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="480" birthdate="2007-01-01" firstname="Jannik" gender="M" lastname="Thiel" license="420091"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="6" heatid="75" lane="3" points="386" resultid="561" swimtime="00:01:07.90"><SPLITS><SPLIT distance="50" swimtime="00:00:31.29"/></SPLITS></RESULT><RESULT eventid="10" heatid="152" lane="2" points="446" resultid="1147" swimtime="00:00:27.35"><SPLITS/></RESULT><RESULT eventid="12" heatid="187" lane="8" points="373" resultid="1419" swimtime="00:02:38.30"><SPLITS><SPLIT distance="50" swimtime="00:00:31.32"/><SPLIT distance="100" swimtime="00:01:13.06"/><SPLIT distance="150" swimtime="00:02:04.32"/></SPLITS></RESULT><RESULT eventid="28" heatid="285" lane="8" points="354" resultid="2123" swimtime="00:00:33.49"><SPLITS/></RESULT><RESULT eventid="30" heatid="322" lane="2" points="429" resultid="2397" swimtime="00:02:15.24"><SPLITS><SPLIT distance="50" swimtime="00:00:31.54"/><SPLIT distance="100" swimtime="00:01:06.53"/><SPLIT distance="150" swimtime="00:01:41.67"/></SPLITS></RESULT><RESULT eventid="36" heatid="396" lane="5" points="477" resultid="2954" swimtime="00:00:28.49"><SPLITS/></RESULT><RESULT eventid="40" heatid="470" lane="6" points="485" resultid="3519" swimtime="00:00:59.62"><SPLITS><SPLIT distance="50" swimtime="00:00:28.95"/></SPLITS></RESULT></RESULTS></ATHLETE></ATHLETES><RELAYS/></CLUB><CLUB code="4360" name="SV Lohhof" nation="GER" region="02" shortname="Lohhof" type="CLUB"><CONTACT city="Unterschleißheim" country="GER" email="johannesbick@hotmail.de" name="Bick, Johannes" street="Carl-von-Linde-Str. 5" zip="85716"/><OFFICIALS/><ATHLETES><ATHLETE athleteid="34" birthdate="2014-01-01" firstname="Anna" gender="F" lastname="Hochstatter" license="460367"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="5" lane="6" points="150" resultid="34" swimtime="00:00:55.09"><SPLITS/></RESULT><RESULT eventid="9" heatid="107" lane="7" points="151" resultid="807" swimtime="00:00:44.43"><SPLITS/></RESULT><RESULT eventid="11" heatid="158" lane="6" points="116" resultid="1195" swimtime="00:04:18.49"><SPLITS><SPLIT distance="50" swimtime="00:01:06.26"/><SPLIT distance="100" swimtime="00:02:10.11"/><SPLIT distance="150" swimtime="00:03:19.68"/></SPLITS></RESULT><RESULT eventid="13" heatid="191" lane="5" points="132" resultid="1444" swimtime="00:01:52.76"><SPLITS><SPLIT distance="50" swimtime="00:00:55.35"/></SPLITS></RESULT><RESULT eventid="21" heatid="237" lane="3" resultid="1776" swimtime="00:01:37.29"><SPLITS/></RESULT><RESULT eventid="23" heatid="240" lane="3" resultid="1790" swimtime="00:01:28.02"><SPLITS/></RESULT><RESULT eventid="31" heatid="328" lane="5" points="136" resultid="2439" swimtime="00:02:04.52"><SPLITS><SPLIT distance="50" swimtime="00:00:56.76"/></SPLITS></RESULT><RESULT eventid="35" heatid="364" lane="2" points="48" resultid="2704" swimtime="00:01:06.88"><SPLITS/></RESULT><RESULT eventid="39" heatid="423" lane="4" points="126" resultid="3150" swimtime="00:01:43.05"><SPLITS><SPLIT distance="50" swimtime="00:00:48.36"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="102" birthdate="2014-01-01" firstname="Pauline" gender="F" lastname="Lettner" license="460369"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="14" lane="2" points="272" resultid="102" swimtime="00:00:45.17"><SPLITS/></RESULT><RESULT eventid="3" heatid="46" lane="6" points="336" resultid="349" swimtime="00:05:39.75"><SPLITS><SPLIT distance="100" swimtime="00:01:22.40"/><SPLIT distance="200" swimtime="00:02:49.78"/><SPLIT distance="300" swimtime="00:04:17.03"/></SPLITS></RESULT><RESULT eventid="7" heatid="85" lane="1" points="232" resultid="633" swimtime="00:03:45.92"><SPLITS><SPLIT distance="50" swimtime="00:00:54.10"/><SPLIT distance="100" swimtime="00:01:49.67"/><SPLIT distance="150" swimtime="00:02:49.49"/></SPLITS></RESULT><RESULT eventid="9" heatid="115" lane="6" points="296" resultid="870" swimtime="00:00:35.50"><SPLITS/></RESULT><RESULT eventid="11" heatid="163" lane="8" points="259" resultid="1234" swimtime="00:03:17.78"><SPLITS><SPLIT distance="50" swimtime="00:00:47.73"/><SPLIT distance="100" swimtime="00:01:39.36"/><SPLIT distance="150" swimtime="00:02:35.87"/></SPLITS></RESULT><RESULT eventid="19" heatid="235" lane="1" resultid="1762" swimtime="00:01:08.05"><SPLITS/></RESULT><RESULT eventid="25" heatid="249" lane="5" resultid="1849" swimtime="00:01:01.28"><SPLITS/></RESULT><RESULT eventid="29" heatid="298" lane="7" points="349" resultid="2220" swimtime="00:02:40.33"><SPLITS><SPLIT distance="50" swimtime="00:00:37.64"/><SPLIT distance="100" swimtime="00:01:19.41"/><SPLIT distance="150" swimtime="00:02:00.58"/></SPLITS></RESULT><RESULT eventid="31" heatid="335" lane="1" points="233" resultid="2491" swimtime="00:01:44.10"><SPLITS><SPLIT distance="50" swimtime="00:00:49.97"/></SPLITS></RESULT><RESULT eventid="35" heatid="366" lane="5" points="204" resultid="2723" swimtime="00:00:41.47"><SPLITS/></RESULT><RESULT eventid="39" heatid="434" lane="4" points="269" resultid="3237" swimtime="00:01:20.03"><SPLITS><SPLIT distance="50" swimtime="00:00:38.37"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="119" birthdate="2010-01-01" firstname="Louisa" gender="F" lastname="Seeber" license="418040"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="16" lane="3" points="222" resultid="119" swimtime="00:00:48.32"><SPLITS/></RESULT><RESULT eventid="3" heatid="41" lane="7" points="233" resultid="311" swimtime="00:06:23.83"><SPLITS><SPLIT distance="200" swimtime="00:03:07.08"/><SPLIT distance="300" swimtime="00:04:46.37"/></SPLITS></RESULT><RESULT eventid="9" heatid="115" lane="7" points="284" resultid="871" swimtime="00:00:36.00"><SPLITS/></RESULT><RESULT eventid="11" heatid="162" lane="1" points="219" resultid="1219" swimtime="00:03:29.22"><SPLITS><SPLIT distance="50" swimtime="00:00:44.44"/><SPLIT distance="100" swimtime="00:01:40.63"/><SPLIT distance="150" swimtime="00:02:41.91"/></SPLITS></RESULT><RESULT eventid="13" heatid="199" lane="1" points="236" resultid="1504" swimtime="00:01:32.93"><SPLITS><SPLIT distance="50" swimtime="00:00:45.78"/></SPLITS></RESULT><RESULT eventid="29" heatid="292" lane="7" points="256" resultid="2172" swimtime="00:02:57.92"><SPLITS><SPLIT distance="50" swimtime="00:00:39.27"/><SPLIT distance="100" swimtime="00:01:25.23"/><SPLIT distance="150" swimtime="00:02:11.51"/></SPLITS></RESULT><RESULT eventid="31" heatid="337" lane="4" points="233" resultid="2510" swimtime="00:01:44.12"><SPLITS><SPLIT distance="50" swimtime="00:00:49.69"/></SPLITS></RESULT><RESULT eventid="35" heatid="370" lane="6" points="204" resultid="2756" swimtime="00:00:41.47"><SPLITS/></RESULT><RESULT eventid="39" heatid="432" lane="6" points="230" resultid="3223" swimtime="00:01:24.37"><SPLITS><SPLIT distance="50" swimtime="00:00:39.56"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="126" birthdate="2011-01-01" firstname="Amelie" gender="F" lastname="Buckl" license="429640"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="17" lane="2" points="292" resultid="126" swimtime="00:00:44.12"><SPLITS/></RESULT><RESULT eventid="5" heatid="65" lane="8" points="147" resultid="488" swimtime="00:01:45.05"><SPLITS><SPLIT distance="50" swimtime="00:00:46.02"/></SPLITS></RESULT><RESULT eventid="7" heatid="88" lane="7" points="287" resultid="663" swimtime="00:03:30.55"><SPLITS><SPLIT distance="50" swimtime="00:00:47.52"/><SPLIT distance="100" swimtime="00:01:41.75"/><SPLIT distance="150" swimtime="00:02:38.03"/></SPLITS></RESULT><RESULT eventid="9" heatid="116" lane="2" points="310" resultid="874" swimtime="00:00:34.97"><SPLITS/></RESULT><RESULT eventid="11" heatid="162" lane="6" points="282" resultid="1224" swimtime="00:03:12.30"><SPLITS><SPLIT distance="50" swimtime="00:00:42.47"/><SPLIT distance="100" swimtime="00:01:32.67"/><SPLIT distance="150" swimtime="00:02:28.49"/></SPLITS></RESULT><RESULT eventid="17" heatid="230" lane="8" points="260" resultid="1739" swimtime="00:12:39.12"><SPLITS><SPLIT distance="100" swimtime="00:01:25.18"/><SPLIT distance="200" swimtime="00:02:59.53"/><SPLIT distance="300" swimtime="00:04:36.19"/><SPLIT distance="400" swimtime="00:06:12.43"/><SPLIT distance="500" swimtime="00:07:50.92"/><SPLIT distance="600" swimtime="00:09:29.16"/><SPLIT distance="700" swimtime="00:11:05.88"/></SPLITS></RESULT><RESULT eventid="27" heatid="264" lane="7" points="291" resultid="1962" swimtime="00:00:40.69"><SPLITS/></RESULT><RESULT eventid="31" heatid="337" lane="2" points="277" resultid="2508" swimtime="00:01:38.32"><SPLITS><SPLIT distance="50" swimtime="00:00:46.88"/></SPLITS></RESULT><RESULT eventid="35" heatid="371" lane="2" points="211" resultid="2760" swimtime="00:00:40.99"><SPLITS/></RESULT><RESULT eventid="39" heatid="434" lane="7" points="307" resultid="3240" swimtime="00:01:16.60"><SPLITS><SPLIT distance="50" swimtime="00:00:36.26"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="136" birthdate="2009-01-01" firstname="Emma" gender="F" lastname="Laux" license="374333"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="18" lane="4" points="323" resultid="136" swimtime="00:00:42.70"><SPLITS/></RESULT><RESULT eventid="3" heatid="47" lane="2" points="367" resultid="353" swimtime="00:05:30.10"><SPLITS><SPLIT distance="100" swimtime="00:01:15.52"/><SPLIT distance="200" swimtime="00:02:41.31"/><SPLIT distance="300" swimtime="00:04:08.20"/></SPLITS></RESULT><RESULT eventid="5" heatid="67" lane="4" points="291" resultid="499" swimtime="00:01:23.68"><SPLITS><SPLIT distance="50" swimtime="00:00:36.71"/></SPLITS></RESULT><RESULT eventid="9" heatid="127" lane="7" points="450" resultid="965" swimtime="00:00:30.88"><SPLITS/></RESULT><RESULT eventid="11" heatid="169" lane="7" points="357" resultid="1281" swimtime="00:02:57.78"><SPLITS><SPLIT distance="50" swimtime="00:00:39.21"/><SPLIT distance="100" swimtime="00:01:25.38"/><SPLIT distance="150" swimtime="00:02:19.10"/></SPLITS></RESULT><RESULT eventid="27" heatid="266" lane="3" points="313" resultid="1974" swimtime="00:00:39.71"><SPLITS/></RESULT><RESULT eventid="29" heatid="302" lane="2" points="395" resultid="2246" swimtime="00:02:33.91"><SPLITS><SPLIT distance="50" swimtime="00:00:34.32"/><SPLIT distance="100" swimtime="00:01:13.38"/><SPLIT distance="150" swimtime="00:01:55.29"/></SPLITS></RESULT><RESULT eventid="35" heatid="376" lane="3" points="338" resultid="2800" swimtime="00:00:35.05"><SPLITS/></RESULT><RESULT eventid="39" heatid="446" lane="2" points="419" resultid="3329" swimtime="00:01:09.07"><SPLITS><SPLIT distance="50" swimtime="00:00:33.03"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="139" birthdate="2006-01-01" firstname="Lea" gender="F" lastname="Wommelsdorf" license="369803"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="18" lane="7" points="286" resultid="139" swimtime="00:00:44.43"><SPLITS/></RESULT><RESULT eventid="5" heatid="66" lane="4" points="283" resultid="492" swimtime="00:01:24.47"><SPLITS><SPLIT distance="50" swimtime="00:00:37.51"/></SPLITS></RESULT><RESULT eventid="11" heatid="168" lane="4" points="347" resultid="1270" swimtime="00:02:59.44"><SPLITS><SPLIT distance="50" swimtime="00:00:36.20"/><SPLIT distance="100" swimtime="00:01:21.67"/><SPLIT distance="150" swimtime="00:02:17.12"/></SPLITS></RESULT><RESULT eventid="13" heatid="207" lane="8" points="369" resultid="1574" swimtime="00:01:20.07"><SPLITS><SPLIT distance="50" swimtime="00:00:38.69"/></SPLITS></RESULT><RESULT eventid="17" heatid="230" lane="3" points="348" resultid="1734" swimtime="00:11:28.66"><SPLITS><SPLIT distance="100" swimtime="00:01:14.44"/><SPLIT distance="200" swimtime="00:02:39.65"/><SPLIT distance="300" swimtime="00:04:06.95"/><SPLIT distance="400" swimtime="00:05:35.92"/><SPLIT distance="500" swimtime="00:07:05.07"/><SPLIT distance="600" swimtime="00:08:34.34"/><SPLIT distance="700" swimtime="00:10:02.67"/></SPLITS></RESULT><RESULT eventid="27" heatid="268" lane="4" points="383" resultid="1991" swimtime="00:00:37.12"><SPLITS/></RESULT><RESULT eventid="31" heatid="339" lane="1" points="271" resultid="2523" swimtime="00:01:39.07"><SPLITS><SPLIT distance="50" swimtime="00:00:47.74"/></SPLITS></RESULT><RESULT eventid="37" heatid="408" lane="5" points="357" resultid="3043" swimtime="00:02:53.85"><SPLITS><SPLIT distance="50" swimtime="00:00:40.36"/><SPLIT distance="100" swimtime="00:01:24.12"/><SPLIT distance="150" swimtime="00:02:10.80"/></SPLITS></RESULT><RESULT eventid="39" heatid="442" lane="4" points="324" resultid="3300" swimtime="00:01:15.23"><SPLITS><SPLIT distance="50" swimtime="00:00:34.75"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="184" birthdate="2010-01-01" firstname="Fiona" gender="F" lastname="Kuhn" license="456503"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="24" lane="6" points="473" resultid="184" swimtime="00:00:37.60"><SPLITS/></RESULT><RESULT eventid="5" heatid="66" lane="7" points="330" resultid="495" swimtime="00:01:20.24"><SPLITS><SPLIT distance="50" swimtime="00:00:36.19"/></SPLITS></RESULT><RESULT eventid="7" heatid="91" lane="2" points="389" resultid="682" swimtime="00:03:10.28"><SPLITS><SPLIT distance="50" swimtime="00:00:41.46"/><SPLIT distance="100" swimtime="00:01:27.80"/><SPLIT distance="150" swimtime="00:02:19.70"/></SPLITS></RESULT><RESULT eventid="9" heatid="126" lane="4" points="449" resultid="955" swimtime="00:00:30.90"><SPLITS/></RESULT><RESULT eventid="11" heatid="168" lane="3" points="402" resultid="1269" swimtime="00:02:50.81"><SPLITS><SPLIT distance="50" swimtime="00:00:36.77"/><SPLIT distance="100" swimtime="00:01:23.18"/><SPLIT distance="150" swimtime="00:02:11.27"/></SPLITS></RESULT><RESULT eventid="17" heatid="230" lane="1" points="337" resultid="1732" swimtime="00:11:36.06"><SPLITS><SPLIT distance="100" swimtime="00:01:15.85"/><SPLIT distance="200" swimtime="00:02:43.19"/><SPLIT distance="300" swimtime="00:04:11.84"/><SPLIT distance="400" swimtime="00:05:41.94"/><SPLIT distance="500" swimtime="00:07:12.96"/><SPLIT distance="600" swimtime="00:08:43.57"/><SPLIT distance="700" swimtime="00:10:11.43"/></SPLITS></RESULT><RESULT eventid="27" heatid="267" lane="6" points="379" resultid="1985" swimtime="00:00:37.25"><SPLITS/></RESULT><RESULT eventid="29" heatid="300" lane="2" points="391" resultid="2231" swimtime="00:02:34.48"><SPLITS><SPLIT distance="50" swimtime="00:00:35.19"/><SPLIT distance="100" swimtime="00:01:14.13"/><SPLIT distance="150" swimtime="00:01:55.10"/></SPLITS></RESULT><RESULT eventid="31" heatid="343" lane="5" points="415" resultid="2559" swimtime="00:01:25.93"><SPLITS><SPLIT distance="50" swimtime="00:00:39.25"/></SPLITS></RESULT><RESULT eventid="35" heatid="373" lane="1" points="320" resultid="2775" swimtime="00:00:35.71"><SPLITS/></RESULT><RESULT eventid="39" heatid="441" lane="5" points="410" resultid="3293" swimtime="00:01:09.58"><SPLITS><SPLIT distance="50" swimtime="00:00:33.40"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="242" birthdate="2014-01-01" firstname="Jan" gender="M" lastname="Brkic" license="460366"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="32" lane="6" points="161" resultid="242" swimtime="00:00:47.63"><SPLITS/></RESULT><RESULT eventid="6" heatid="72" lane="8" points="107" resultid="543" swimtime="00:01:43.88"><SPLITS><SPLIT distance="50" swimtime="00:00:45.34"/></SPLITS></RESULT><RESULT eventid="8" heatid="95" lane="6" points="174" resultid="715" swimtime="00:03:45.21"><SPLITS><SPLIT distance="50" swimtime="00:00:52.13"/><SPLIT distance="100" swimtime="00:01:49.11"/><SPLIT distance="150" swimtime="00:02:47.31"/></SPLITS></RESULT><RESULT eventid="10" heatid="143" lane="8" points="244" resultid="1081" swimtime="00:00:33.46"><SPLITS/></RESULT><RESULT eventid="14" heatid="217" lane="4" points="188" resultid="1646" swimtime="00:01:29.94"><SPLITS><SPLIT distance="50" swimtime="00:00:42.66"/></SPLITS></RESULT><RESULT eventid="18" heatid="232" lane="6" points="295" resultid="1752" swimtime="00:11:18.68"><SPLITS><SPLIT distance="100" swimtime="00:01:19.73"/><SPLIT distance="200" swimtime="00:02:45.48"/><SPLIT distance="300" swimtime="00:04:12.15"/><SPLIT distance="400" swimtime="00:05:39.93"/><SPLIT distance="500" swimtime="00:07:06.26"/><SPLIT distance="600" swimtime="00:08:32.97"/><SPLIT distance="700" swimtime="00:09:59.14"/></SPLITS></RESULT><RESULT eventid="22" heatid="239" lane="5" resultid="1788" swimtime="00:01:00.69"><SPLITS/></RESULT><RESULT comment="08:52 Start vor dem Startsignal" eventid="24" heatid="245" lane="3" resultid="1822" status="DSQ" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="26" heatid="251" lane="6" resultid="1860" swimtime="00:00:59.44"><SPLITS/></RESULT><RESULT eventid="32" heatid="349" lane="4" points="158" resultid="2600" swimtime="00:01:45.06"><SPLITS><SPLIT distance="50" swimtime="00:00:50.23"/></SPLITS></RESULT><RESULT eventid="36" heatid="387" lane="8" points="127" resultid="2885" swimtime="00:00:44.19"><SPLITS/></RESULT><RESULT eventid="40" heatid="462" lane="8" points="254" resultid="3459" swimtime="00:01:13.94"><SPLITS><SPLIT distance="50" swimtime="00:00:35.91"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="394" birthdate="2013-01-01" firstname="Domenik" gender="M" lastname="Pavlitschek" license="457421"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="56" lane="1" points="229" resultid="418" swimtime="00:05:59.31"><SPLITS><SPLIT distance="100" swimtime="00:01:25.03"/><SPLIT distance="200" swimtime="00:02:56.50"/><SPLIT distance="300" swimtime="00:04:28.09"/></SPLITS></RESULT><RESULT eventid="6" heatid="72" lane="5" points="111" resultid="540" swimtime="00:01:42.59"><SPLITS><SPLIT distance="50" swimtime="00:00:44.86"/></SPLITS></RESULT><RESULT eventid="10" heatid="142" lane="3" points="198" resultid="1069" swimtime="00:00:35.83"><SPLITS/></RESULT><RESULT eventid="12" heatid="178" lane="8" points="190" resultid="1349" swimtime="00:03:18.00"><SPLITS><SPLIT distance="50" swimtime="00:00:47.89"/><SPLIT distance="100" swimtime="00:01:39.22"/><SPLIT distance="150" swimtime="00:02:36.47"/></SPLITS></RESULT><RESULT eventid="14" heatid="216" lane="6" points="156" resultid="1640" swimtime="00:01:35.84"><SPLITS><SPLIT distance="50" swimtime="00:00:46.68"/></SPLITS></RESULT><RESULT eventid="22" heatid="239" lane="3" resultid="1786" swimtime="00:01:07.01"><SPLITS/></RESULT><RESULT eventid="24" heatid="244" lane="4" resultid="1817" swimtime="00:00:55.37"><SPLITS/></RESULT><RESULT comment="09:07 Der Sportler führte nach dem Start mehrere Wechselbeinschläge durch" eventid="26" heatid="251" lane="4" resultid="1858" status="DSQ" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="32" heatid="349" lane="8" points="144" resultid="2604" swimtime="00:01:48.27"><SPLITS><SPLIT distance="50" swimtime="00:00:52.32"/></SPLITS></RESULT><RESULT eventid="36" heatid="385" lane="5" points="149" resultid="2867" swimtime="00:00:41.98"><SPLITS/></RESULT><RESULT eventid="40" heatid="460" lane="6" points="206" resultid="3441" swimtime="00:01:19.34"><SPLITS><SPLIT distance="50" swimtime="00:00:37.81"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="418" birthdate="2010-01-01" firstname="Tim Julius" gender="M" lastname="Listing" license="441345"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="59" lane="7" points="328" resultid="447" swimtime="00:05:19.02"><SPLITS><SPLIT distance="100" swimtime="00:01:10.62"/><SPLIT distance="200" swimtime="00:02:32.80"/><SPLIT distance="300" swimtime="00:03:57.20"/></SPLITS></RESULT><RESULT eventid="6" heatid="75" lane="6" points="239" resultid="564" swimtime="00:01:19.61"><SPLITS><SPLIT distance="50" swimtime="00:00:34.80"/></SPLITS></RESULT><RESULT eventid="10" heatid="148" lane="8" points="372" resultid="1121" swimtime="00:00:29.05"><SPLITS/></RESULT><RESULT eventid="12" heatid="185" lane="1" points="329" resultid="1396" swimtime="00:02:45.11"><SPLITS><SPLIT distance="50" swimtime="00:00:35.41"/><SPLIT distance="100" swimtime="00:01:17.93"/><SPLIT distance="150" swimtime="00:02:09.67"/></SPLITS></RESULT><RESULT eventid="14" heatid="222" lane="1" points="306" resultid="1682" swimtime="00:01:16.51"><SPLITS><SPLIT distance="50" swimtime="00:00:37.87"/></SPLITS></RESULT><RESULT eventid="28" heatid="284" lane="1" points="293" resultid="2109" swimtime="00:00:35.69"><SPLITS/></RESULT><RESULT eventid="30" heatid="321" lane="5" points="369" resultid="2392" swimtime="00:02:22.19"><SPLITS><SPLIT distance="50" swimtime="00:00:31.05"/><SPLIT distance="100" swimtime="00:01:06.89"/><SPLIT distance="150" swimtime="00:01:45.41"/></SPLITS></RESULT><RESULT eventid="36" heatid="393" lane="1" points="301" resultid="2926" swimtime="00:00:33.21"><SPLITS/></RESULT><RESULT eventid="40" heatid="468" lane="5" points="394" resultid="3502" swimtime="00:01:03.91"><SPLITS><SPLIT distance="50" swimtime="00:00:30.92"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="440" birthdate="2013-01-01" firstname="Lina" gender="F" lastname="Janotta" license="456507"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="5" heatid="64" lane="1" points="139" resultid="473" swimtime="00:01:46.95"><SPLITS><SPLIT distance="50" swimtime="00:00:46.29"/></SPLITS></RESULT><RESULT eventid="9" heatid="118" lane="2" points="421" resultid="889" swimtime="00:00:31.57"><SPLITS/></RESULT><RESULT eventid="11" heatid="161" lane="2" points="308" resultid="1212" swimtime="00:03:06.65"><SPLITS><SPLIT distance="50" swimtime="00:00:40.33"/><SPLIT distance="100" swimtime="00:01:25.46"/><SPLIT distance="150" swimtime="00:02:25.85"/></SPLITS></RESULT><RESULT eventid="13" heatid="204" lane="1" points="327" resultid="1544" swimtime="00:01:23.36"><SPLITS><SPLIT distance="50" swimtime="00:00:40.10"/></SPLITS></RESULT><RESULT eventid="17" heatid="230" lane="7" resultid="1738" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="19" heatid="235" lane="5" resultid="1766" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="21" heatid="238" lane="4" resultid="1781" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="23" heatid="243" lane="1" resultid="1807" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="29" heatid="298" lane="6" resultid="2219" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="37" heatid="408" lane="1" resultid="3039" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="39" heatid="437" lane="2" resultid="3259" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="532" birthdate="2004-01-01" firstname="Evelin" gender="F" lastname="Laux" license="334210"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="9" heatid="129" lane="8" points="476" resultid="982" swimtime="00:00:30.30"><SPLITS/></RESULT><RESULT eventid="35" heatid="380" lane="7" points="380" resultid="2834" swimtime="00:00:33.70"><SPLITS/></RESULT></RESULTS></ATHLETE></ATHLETES><RELAYS/></CLUB><CLUB code="6524" name="SC Regensburg" nation="GER" region="02" shortname="Regensbg" type="CLUB"><CONTACT city="Regensburg" country="GER" email="julia.bauer@sc-rgbg.de" name="Bauer, Julia" phone="0941/37805208" street="Messerschmittstr. 4" zip="93049"/><OFFICIALS/><ATHLETES><ATHLETE athleteid="35" birthdate="2014-01-01" firstname="Charlotte" gender="F" lastname="Walz" license="449243"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="5" lane="7" points="144" resultid="35" swimtime="00:00:55.87"><SPLITS/></RESULT><RESULT eventid="9" heatid="108" lane="2" points="120" resultid="810" swimtime="00:00:47.92"><SPLITS/></RESULT><RESULT eventid="13" heatid="191" lane="4" points="122" resultid="1443" swimtime="00:01:55.68"><SPLITS/></RESULT><RESULT eventid="29" heatid="290" lane="6" points="135" resultid="2156" swimtime="00:03:39.73"><SPLITS><SPLIT distance="50" swimtime="00:00:46.34"/><SPLIT distance="100" swimtime="00:01:43.21"/><SPLIT distance="150" swimtime="00:02:43.69"/></SPLITS></RESULT><RESULT eventid="35" heatid="363" lane="7" points="77" resultid="2701" swimtime="00:00:57.18"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="38" birthdate="2016-01-01" firstname="Leonie" gender="F" lastname="Gierl" license="482482"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="6" lane="2" points="123" resultid="38" swimtime="00:00:58.76"><SPLITS/></RESULT><RESULT eventid="9" heatid="103" lane="7" points="92" resultid="775" swimtime="00:00:52.34"><SPLITS/></RESULT><RESULT eventid="13" heatid="190" lane="6" points="103" resultid="1439" swimtime="00:02:02.39"><SPLITS><SPLIT distance="50" swimtime="00:00:57.28"/></SPLITS></RESULT><RESULT eventid="27" heatid="253" lane="4" points="118" resultid="1871" swimtime="00:00:54.99"><SPLITS/></RESULT><RESULT eventid="31" heatid="328" lane="6" points="131" resultid="2440" swimtime="00:02:06.05"><SPLITS><SPLIT distance="50" swimtime="00:00:59.38"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="39" birthdate="2014-01-01" firstname="Louisa" gender="F" lastname="Muñoz" license="457808"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="6" lane="3" points="173" resultid="39" swimtime="00:00:52.51"><SPLITS/></RESULT><RESULT eventid="7" heatid="82" lane="3" points="203" resultid="612" swimtime="00:03:56.09"><SPLITS><SPLIT distance="50" swimtime="00:00:54.13"/><SPLIT distance="100" swimtime="00:01:54.16"/><SPLIT distance="150" swimtime="00:02:57.18"/></SPLITS></RESULT><RESULT eventid="9" heatid="111" lane="8" points="220" resultid="840" swimtime="00:00:39.19"><SPLITS/></RESULT><RESULT eventid="13" heatid="198" lane="1" points="217" resultid="1496" swimtime="00:01:35.56"><SPLITS><SPLIT distance="50" swimtime="00:00:48.36"/></SPLITS></RESULT><RESULT eventid="29" heatid="294" lane="7" points="239" resultid="2188" swimtime="00:03:01.86"><SPLITS><SPLIT distance="50" swimtime="00:00:40.93"/><SPLIT distance="100" swimtime="00:01:29.06"/><SPLIT distance="150" swimtime="00:02:17.09"/></SPLITS></RESULT><RESULT eventid="31" heatid="333" lane="4" points="178" resultid="2478" swimtime="00:01:53.92"><SPLITS><SPLIT distance="50" swimtime="00:00:53.86"/></SPLITS></RESULT><RESULT eventid="35" heatid="368" lane="6" points="185" resultid="2740" swimtime="00:00:42.84"><SPLITS/></RESULT><RESULT eventid="39" heatid="431" lane="8" points="228" resultid="3217" swimtime="00:01:24.64"><SPLITS><SPLIT distance="50" swimtime="00:00:41.86"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="40" birthdate="2015-01-01" firstname="Sofía" gender="F" lastname="Hutchinson Riquelme" license="472000"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="6" lane="4" points="144" resultid="40" swimtime="00:00:55.81"><SPLITS/></RESULT><RESULT eventid="7" heatid="81" lane="2" points="171" resultid="605" swimtime="00:04:09.92"><SPLITS><SPLIT distance="50" swimtime="00:00:57.91"/><SPLIT distance="100" swimtime="00:02:00.67"/><SPLIT distance="150" swimtime="00:03:05.97"/></SPLITS></RESULT><RESULT eventid="9" heatid="105" lane="3" points="105" resultid="787" swimtime="00:00:50.03"><SPLITS/></RESULT><RESULT eventid="13" heatid="192" lane="7" points="103" resultid="1454" swimtime="00:02:02.44"><SPLITS><SPLIT distance="50" swimtime="00:01:01.22"/></SPLITS></RESULT><RESULT eventid="27" heatid="256" lane="1" points="115" resultid="1892" swimtime="00:00:55.37"><SPLITS/></RESULT><RESULT eventid="31" heatid="329" lane="5" points="154" resultid="2447" swimtime="00:01:59.45"><SPLITS><SPLIT distance="50" swimtime="00:00:57.31"/></SPLITS></RESULT><RESULT eventid="39" heatid="422" lane="5" points="109" resultid="3143" swimtime="00:01:48.22"><SPLITS><SPLIT distance="50" swimtime="00:00:50.80"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="63" birthdate="2014-01-01" firstname="Lucy" gender="F" lastname="Song" license="449372"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="9" lane="3" points="150" resultid="63" swimtime="00:00:55.09"><SPLITS/></RESULT><RESULT eventid="13" heatid="193" lane="1" points="163" resultid="1456" swimtime="00:01:45.04"><SPLITS><SPLIT distance="50" swimtime="00:00:50.26"/></SPLITS></RESULT><RESULT eventid="27" heatid="259" lane="4" points="160" resultid="1919" swimtime="00:00:49.63"><SPLITS/></RESULT><RESULT eventid="29" heatid="288" lane="2" points="108" resultid="2138" swimtime="00:03:56.65"><SPLITS><SPLIT distance="50" swimtime="00:00:48.00"/><SPLIT distance="100" swimtime="00:01:48.13"/><SPLIT distance="150" swimtime="00:02:53.26"/></SPLITS></RESULT><RESULT eventid="31" heatid="329" lane="7" points="155" resultid="2449" swimtime="00:01:59.22"><SPLITS><SPLIT distance="50" swimtime="00:00:55.42"/></SPLITS></RESULT><RESULT eventid="39" heatid="423" lane="8" points="134" resultid="3154" swimtime="00:01:41.00"><SPLITS><SPLIT distance="50" swimtime="00:00:47.08"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="72" birthdate="2015-01-01" firstname="Anna" gender="F" lastname="Stendel" license="464758"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="10" lane="4" points="207" resultid="72" swimtime="00:00:49.47"><SPLITS/></RESULT><RESULT eventid="7" heatid="82" lane="5" points="193" resultid="614" swimtime="00:04:00.05"><SPLITS><SPLIT distance="50" swimtime="00:00:52.49"/><SPLIT distance="100" swimtime="00:01:54.01"/><SPLIT distance="150" swimtime="00:02:58.09"/></SPLITS></RESULT><RESULT eventid="9" heatid="110" lane="6" points="196" resultid="830" swimtime="00:00:40.74"><SPLITS/></RESULT><RESULT eventid="13" heatid="194" lane="8" points="149" resultid="1471" swimtime="00:01:48.18"><SPLITS><SPLIT distance="50" swimtime="00:00:54.63"/></SPLITS></RESULT><RESULT eventid="27" heatid="258" lane="6" points="159" resultid="1913" swimtime="00:00:49.78"><SPLITS/></RESULT><RESULT eventid="31" heatid="332" lane="5" points="189" resultid="2471" swimtime="00:01:51.74"><SPLITS><SPLIT distance="50" swimtime="00:00:52.30"/></SPLITS></RESULT><RESULT eventid="35" heatid="363" lane="8" points="70" resultid="2702" swimtime="00:00:59.02"><SPLITS/></RESULT><RESULT eventid="39" heatid="427" lane="6" points="161" resultid="3183" swimtime="00:01:34.98"><SPLITS><SPLIT distance="50" swimtime="00:00:42.90"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="83" birthdate="2015-01-01" firstname="Hanna" gender="F" lastname="Gierl" license="471997"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="11" lane="7" points="198" resultid="83" swimtime="00:00:50.26"><SPLITS/></RESULT><RESULT eventid="7" heatid="85" lane="3" points="232" resultid="635" swimtime="00:03:45.85"><SPLITS><SPLIT distance="50" swimtime="00:00:52.24"/><SPLIT distance="100" swimtime="00:01:52.09"/><SPLIT distance="150" swimtime="00:02:50.04"/></SPLITS></RESULT><RESULT eventid="9" heatid="105" lane="6" points="105" resultid="790" swimtime="00:00:50.11"><SPLITS/></RESULT><RESULT eventid="13" heatid="192" lane="4" points="107" resultid="1451" swimtime="00:02:00.97"><SPLITS><SPLIT distance="50" swimtime="00:00:57.90"/></SPLITS></RESULT><RESULT eventid="27" heatid="256" lane="2" points="132" resultid="1893" swimtime="00:00:52.90"><SPLITS/></RESULT><RESULT eventid="31" heatid="333" lane="6" points="203" resultid="2480" swimtime="00:01:49.02"><SPLITS><SPLIT distance="50" swimtime="00:00:52.38"/></SPLITS></RESULT><RESULT eventid="37" heatid="401" lane="5" points="136" resultid="2991" swimtime="00:03:59.75"><SPLITS><SPLIT distance="50" swimtime="00:00:54.45"/><SPLIT distance="100" swimtime="00:01:58.48"/><SPLIT distance="150" swimtime="00:02:59.45"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="88" birthdate="2014-01-01" firstname="Julia" gender="F" lastname="Rummel" license="458196"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="12" lane="4" points="252" resultid="88" swimtime="00:00:46.34"><SPLITS/></RESULT><RESULT eventid="7" heatid="87" lane="2" points="296" resultid="650" swimtime="00:03:28.42"><SPLITS><SPLIT distance="50" swimtime="00:00:48.11"/><SPLIT distance="100" swimtime="00:01:40.73"/><SPLIT distance="150" swimtime="00:02:36.01"/></SPLITS></RESULT><RESULT eventid="9" heatid="114" lane="2" points="271" resultid="858" swimtime="00:00:36.56"><SPLITS/></RESULT><RESULT eventid="11" heatid="164" lane="3" points="285" resultid="1237" swimtime="00:03:11.60"><SPLITS><SPLIT distance="50" swimtime="00:00:41.70"/><SPLIT distance="100" swimtime="00:01:33.64"/><SPLIT distance="150" swimtime="00:02:28.03"/></SPLITS></RESULT><RESULT eventid="23" heatid="242" lane="6" resultid="1804" swimtime="00:01:02.38"><SPLITS/></RESULT><RESULT eventid="27" heatid="261" lane="5" points="230" resultid="1936" swimtime="00:00:43.98"><SPLITS/></RESULT><RESULT eventid="29" heatid="297" lane="7" points="284" resultid="2212" swimtime="00:02:51.70"><SPLITS><SPLIT distance="50" swimtime="00:00:38.18"/><SPLIT distance="100" swimtime="00:01:22.20"/><SPLIT distance="150" swimtime="00:02:06.80"/></SPLITS></RESULT><RESULT eventid="35" heatid="368" lane="1" points="202" resultid="2735" swimtime="00:00:41.59"><SPLITS/></RESULT><RESULT eventid="39" heatid="432" lane="3" points="263" resultid="3220" swimtime="00:01:20.66"><SPLITS><SPLIT distance="50" swimtime="00:00:38.91"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="91" birthdate="2015-01-01" firstname="Emilia" gender="F" lastname="Soric" license="471993"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="12" lane="7" points="218" resultid="91" swimtime="00:00:48.62"><SPLITS/></RESULT><RESULT eventid="7" heatid="84" lane="1" points="233" resultid="625" swimtime="00:03:45.80"><SPLITS><SPLIT distance="50" swimtime="00:00:53.80"/><SPLIT distance="100" swimtime="00:01:48.92"/><SPLIT distance="150" swimtime="00:02:50.90"/></SPLITS></RESULT><RESULT eventid="9" heatid="107" lane="2" points="127" resultid="802" swimtime="00:00:47.04"><SPLITS/></RESULT><RESULT eventid="27" heatid="253" lane="6" points="180" resultid="1873" swimtime="00:00:47.73"><SPLITS/></RESULT><RESULT eventid="31" heatid="334" lane="2" points="213" resultid="2484" swimtime="00:01:47.36"><SPLITS><SPLIT distance="50" swimtime="00:00:51.77"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="132" birthdate="2012-01-01" firstname="Sophia" gender="F" lastname="Löw" license="442814"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="17" lane="8" points="291" resultid="132" swimtime="00:00:44.21"><SPLITS/></RESULT><RESULT eventid="7" heatid="89" lane="8" points="333" resultid="672" swimtime="00:03:20.41"><SPLITS><SPLIT distance="50" swimtime="00:00:47.79"/><SPLIT distance="100" swimtime="00:01:39.26"/><SPLIT distance="150" swimtime="00:02:31.66"/></SPLITS></RESULT><RESULT eventid="9" heatid="117" lane="1" points="328" resultid="881" swimtime="00:00:34.31"><SPLITS/></RESULT><RESULT eventid="13" heatid="197" lane="7" points="239" resultid="1494" swimtime="00:01:32.56"><SPLITS><SPLIT distance="50" swimtime="00:00:45.29"/></SPLITS></RESULT><RESULT eventid="29" heatid="298" lane="4" points="349" resultid="2217" swimtime="00:02:40.41"><SPLITS><SPLIT distance="50" swimtime="00:00:37.39"/><SPLIT distance="100" swimtime="00:01:20.18"/><SPLIT distance="150" swimtime="00:02:01.60"/></SPLITS></RESULT><RESULT eventid="31" heatid="338" lane="6" points="312" resultid="2520" swimtime="00:01:34.46"><SPLITS><SPLIT distance="50" swimtime="00:00:45.08"/></SPLITS></RESULT><RESULT eventid="37" heatid="405" lane="3" points="262" resultid="3017" swimtime="00:03:12.71"><SPLITS><SPLIT distance="50" swimtime="00:00:47.80"/><SPLIT distance="100" swimtime="00:01:37.85"/><SPLIT distance="150" swimtime="00:02:27.53"/></SPLITS></RESULT><RESULT eventid="39" heatid="434" lane="2" points="301" resultid="3235" swimtime="00:01:17.14"><SPLITS><SPLIT distance="50" swimtime="00:00:37.35"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="135" birthdate="2011-01-01" firstname="Mia Luisa" gender="F" lastname="Schönberger" license="443832"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="18" lane="3" points="333" resultid="135" swimtime="00:00:42.27"><SPLITS/></RESULT><RESULT eventid="7" heatid="89" lane="3" points="356" resultid="667" swimtime="00:03:16.03"><SPLITS><SPLIT distance="50" swimtime="00:00:45.49"/><SPLIT distance="100" swimtime="00:01:36.03"/><SPLIT distance="150" swimtime="00:02:27.24"/></SPLITS></RESULT><RESULT eventid="13" heatid="206" lane="8" points="392" resultid="1567" swimtime="00:01:18.47"><SPLITS><SPLIT distance="50" swimtime="00:00:37.98"/></SPLITS></RESULT><RESULT eventid="27" heatid="268" lane="3" points="423" resultid="1990" swimtime="00:00:35.93"><SPLITS/></RESULT><RESULT eventid="31" heatid="339" lane="3" points="331" resultid="2525" swimtime="00:01:32.64"><SPLITS><SPLIT distance="50" swimtime="00:00:45.23"/></SPLITS></RESULT><RESULT eventid="37" heatid="408" lane="2" points="373" resultid="3040" swimtime="00:02:51.22"><SPLITS><SPLIT distance="50" swimtime="00:00:38.44"/><SPLIT distance="100" swimtime="00:01:22.56"/><SPLIT distance="150" swimtime="00:02:08.01"/></SPLITS></RESULT><RESULT eventid="39" heatid="438" lane="1" points="378" resultid="3266" swimtime="00:01:11.46"><SPLITS><SPLIT distance="50" swimtime="00:00:34.67"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="148" birthdate="2013-01-01" firstname="Johanna" gender="F" lastname="Spitzner" license="443850"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="19" lane="8" points="326" resultid="148" swimtime="00:00:42.55"><SPLITS/></RESULT><RESULT eventid="7" heatid="84" lane="5" points="325" resultid="629" swimtime="00:03:22.07"><SPLITS><SPLIT distance="50" swimtime="00:00:44.60"/><SPLIT distance="100" swimtime="00:01:38.00"/><SPLIT distance="150" swimtime="00:02:31.18"/></SPLITS></RESULT><RESULT eventid="9" heatid="116" lane="1" points="313" resultid="873" swimtime="00:00:34.83"><SPLITS/></RESULT><RESULT eventid="11" heatid="166" lane="1" points="309" resultid="1251" swimtime="00:03:06.52"><SPLITS><SPLIT distance="50" swimtime="00:00:38.17"/><SPLIT distance="100" swimtime="00:01:29.47"/><SPLIT distance="150" swimtime="00:02:23.68"/></SPLITS></RESULT><RESULT eventid="21" heatid="238" lane="6" resultid="1783" swimtime="00:00:45.51"><SPLITS/></RESULT><RESULT eventid="27" heatid="264" lane="5" points="312" resultid="1960" swimtime="00:00:39.74"><SPLITS/></RESULT><RESULT eventid="29" heatid="296" lane="2" points="255" resultid="2199" swimtime="00:02:58.05"><SPLITS><SPLIT distance="50" swimtime="00:00:38.79"/><SPLIT distance="100" swimtime="00:01:23.27"/><SPLIT distance="150" swimtime="00:02:11.81"/></SPLITS></RESULT><RESULT eventid="37" heatid="406" lane="8" points="289" resultid="3030" swimtime="00:03:06.40"><SPLITS><SPLIT distance="50" swimtime="00:00:44.02"/><SPLIT distance="100" swimtime="00:01:31.18"/><SPLIT distance="150" swimtime="00:02:20.67"/></SPLITS></RESULT><RESULT eventid="39" heatid="436" lane="8" points="294" resultid="3257" swimtime="00:01:17.72"><SPLITS><SPLIT distance="50" swimtime="00:00:37.13"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="150" birthdate="2011-01-01" firstname="Julia Pia" gender="F" lastname="Schüller" license="443830"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="20" lane="2" points="343" resultid="150" swimtime="00:00:41.82"><SPLITS/></RESULT><RESULT eventid="5" heatid="68" lane="6" points="337" resultid="509" swimtime="00:01:19.71"><SPLITS><SPLIT distance="50" swimtime="00:00:35.31"/></SPLITS></RESULT><RESULT eventid="9" heatid="125" lane="5" points="425" resultid="948" swimtime="00:00:31.46"><SPLITS/></RESULT><RESULT eventid="13" heatid="203" lane="4" points="340" resultid="1539" swimtime="00:01:22.26"><SPLITS><SPLIT distance="50" swimtime="00:00:39.23"/></SPLITS></RESULT><RESULT eventid="27" heatid="267" lane="2" points="361" resultid="1981" swimtime="00:00:37.86"><SPLITS/></RESULT><RESULT eventid="35" heatid="379" lane="2" points="362" resultid="2821" swimtime="00:00:34.27"><SPLITS/></RESULT><RESULT eventid="39" heatid="444" lane="3" points="409" resultid="3315" swimtime="00:01:09.64"><SPLITS><SPLIT distance="50" swimtime="00:00:33.49"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="163" birthdate="2010-01-01" firstname="Teresa" gender="F" lastname="Stangelmayer" license="414346"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="21" lane="8" points="382" resultid="163" swimtime="00:00:40.35"><SPLITS/></RESULT><RESULT eventid="7" heatid="91" lane="6" points="474" resultid="686" swimtime="00:02:58.17"><SPLITS><SPLIT distance="50" swimtime="00:00:41.82"/><SPLIT distance="100" swimtime="00:01:26.67"/><SPLIT distance="150" swimtime="00:02:13.15"/></SPLITS></RESULT><RESULT eventid="11" heatid="170" lane="3" points="428" resultid="1285" swimtime="00:02:47.29"><SPLITS><SPLIT distance="50" swimtime="00:00:36.72"/><SPLIT distance="100" swimtime="00:01:23.77"/><SPLIT distance="150" swimtime="00:02:11.31"/></SPLITS></RESULT><RESULT eventid="31" heatid="342" lane="7" points="432" resultid="2553" swimtime="00:01:24.80"><SPLITS><SPLIT distance="50" swimtime="00:00:41.52"/></SPLITS></RESULT><RESULT eventid="35" heatid="378" lane="8" points="363" resultid="2819" swimtime="00:00:34.24"><SPLITS/></RESULT><RESULT eventid="39" heatid="442" lane="7" points="436" resultid="3303" swimtime="00:01:08.15"><SPLITS><SPLIT distance="50" swimtime="00:00:33.08"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="164" birthdate="2012-01-01" firstname="Elisa" gender="F" lastname="Ostermeier" license="442817"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="22" lane="1" points="371" resultid="164" swimtime="00:00:40.76"><SPLITS/></RESULT><RESULT eventid="9" heatid="127" lane="1" points="416" resultid="959" swimtime="00:00:31.69"><SPLITS/></RESULT><RESULT eventid="11" heatid="169" lane="5" points="396" resultid="1279" swimtime="00:02:51.61"><SPLITS><SPLIT distance="50" swimtime="00:00:34.47"/><SPLIT distance="100" swimtime="00:01:20.93"/><SPLIT distance="150" swimtime="00:02:10.67"/></SPLITS></RESULT><RESULT eventid="31" heatid="341" lane="7" points="393" resultid="2545" swimtime="00:01:27.52"><SPLITS><SPLIT distance="50" swimtime="00:00:41.39"/></SPLITS></RESULT><RESULT eventid="35" heatid="375" lane="8" points="331" resultid="2797" swimtime="00:00:35.31"><SPLITS/></RESULT><RESULT eventid="39" heatid="443" lane="8" points="432" resultid="3312" swimtime="00:01:08.38"><SPLITS><SPLIT distance="50" swimtime="00:00:32.61"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="166" birthdate="2009-01-01" firstname="Sarah" gender="F" lastname="Osteroth" license="400513"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="22" lane="3" resultid="166" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="7" heatid="90" lane="8" resultid="680" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="9" heatid="122" lane="4" resultid="923" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="33" heatid="359" lane="1" resultid="2667" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="35" heatid="377" lane="3" resultid="2808" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="174" birthdate="2009-01-01" firstname="Paula" gender="F" lastname="Spitzner" license="400524"><HANDICAP/><ENTRIES/><RESULTS><RESULT comment="09:35 Start vor dem Startsignal" eventid="1" heatid="23" lane="4" resultid="174" status="DSQ" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="7" heatid="92" lane="1" points="464" resultid="689" swimtime="00:02:59.39"><SPLITS><SPLIT distance="50" swimtime="00:00:41.02"/><SPLIT distance="100" swimtime="00:01:25.69"/><SPLIT distance="150" swimtime="00:02:13.29"/></SPLITS></RESULT><RESULT eventid="9" heatid="130" lane="1" points="484" resultid="983" swimtime="00:00:30.13"><SPLITS/></RESULT><RESULT eventid="31" heatid="344" lane="7" points="454" resultid="2569" swimtime="00:01:23.42"><SPLITS><SPLIT distance="50" swimtime="00:00:37.87"/></SPLITS></RESULT><RESULT eventid="35" heatid="380" lane="1" points="369" resultid="2828" swimtime="00:00:34.04"><SPLITS/></RESULT><RESULT eventid="39" heatid="448" lane="4" points="516" resultid="3346" swimtime="00:01:04.43"><SPLITS><SPLIT distance="50" swimtime="00:00:30.28"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="176" birthdate="2011-01-01" firstname="Paula" gender="F" lastname="Rößger" license="442820"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="23" lane="6" points="486" resultid="176" swimtime="00:00:37.25"><SPLITS/></RESULT><RESULT eventid="7" heatid="91" lane="4" points="453" resultid="684" swimtime="00:03:00.80"><SPLITS><SPLIT distance="50" swimtime="00:00:41.32"/><SPLIT distance="100" swimtime="00:01:28.97"/><SPLIT distance="150" swimtime="00:02:15.11"/></SPLITS></RESULT><RESULT eventid="9" heatid="122" lane="3" points="418" resultid="922" swimtime="00:00:31.65"><SPLITS/></RESULT><RESULT eventid="11" heatid="171" lane="7" points="413" resultid="1297" swimtime="00:02:49.22"><SPLITS><SPLIT distance="50" swimtime="00:00:36.80"/><SPLIT distance="100" swimtime="00:01:22.92"/><SPLIT distance="150" swimtime="00:02:11.69"/></SPLITS></RESULT><RESULT eventid="31" heatid="343" lane="3" points="442" resultid="2557" swimtime="00:01:24.16"><SPLITS><SPLIT distance="50" swimtime="00:00:40.83"/></SPLITS></RESULT><RESULT eventid="35" heatid="377" lane="5" points="388" resultid="2809" swimtime="00:00:33.48"><SPLITS/></RESULT><RESULT eventid="39" heatid="445" lane="2" points="435" resultid="3322" swimtime="00:01:08.24"><SPLITS><SPLIT distance="50" swimtime="00:00:32.58"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="201" birthdate="2014-01-01" firstname="Jacob" gender="M" lastname="Mulzer" license="449265"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="27" lane="4" points="130" resultid="201" swimtime="00:00:51.17"><SPLITS/></RESULT><RESULT eventid="8" heatid="94" lane="8" points="151" resultid="711" swimtime="00:03:56.16"><SPLITS><SPLIT distance="50" swimtime="00:00:57.20"/><SPLIT distance="100" swimtime="00:01:57.34"/><SPLIT distance="150" swimtime="00:03:00.74"/></SPLITS></RESULT><RESULT eventid="10" heatid="140" lane="7" points="155" resultid="1058" swimtime="00:00:38.88"><SPLITS/></RESULT><RESULT eventid="14" heatid="215" lane="6" points="140" resultid="1632" swimtime="00:01:39.27"><SPLITS><SPLIT distance="50" swimtime="00:00:47.79"/></SPLITS></RESULT><RESULT eventid="28" heatid="278" lane="3" points="126" resultid="2063" swimtime="00:00:47.22"><SPLITS/></RESULT><RESULT eventid="30" heatid="314" lane="3" points="194" resultid="2336" swimtime="00:02:56.03"><SPLITS><SPLIT distance="50" swimtime="00:00:40.63"/><SPLIT distance="100" swimtime="00:01:25.64"/><SPLIT distance="150" swimtime="00:02:13.09"/></SPLITS></RESULT><RESULT eventid="36" heatid="385" lane="8" points="127" resultid="2870" swimtime="00:00:44.21"><SPLITS/></RESULT><RESULT eventid="40" heatid="459" lane="1" points="165" resultid="3429" swimtime="00:01:25.29"><SPLITS><SPLIT distance="50" swimtime="00:00:40.24"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="205" birthdate="2015-01-01" firstname="Marco" gender="M" lastname="Ivaldi" license="482342"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="28" lane="1" points="108" resultid="205" swimtime="00:00:54.48"><SPLITS/></RESULT><RESULT eventid="10" heatid="135" lane="7" points="87" resultid="1019" swimtime="00:00:47.18"><SPLITS/></RESULT><RESULT eventid="14" heatid="211" lane="5" points="102" resultid="1601" swimtime="00:01:50.40"><SPLITS><SPLIT distance="50" swimtime="00:00:53.84"/></SPLITS></RESULT><RESULT eventid="28" heatid="277" lane="7" points="103" resultid="2059" swimtime="00:00:50.56"><SPLITS/></RESULT><RESULT eventid="30" heatid="308" lane="2" points="83" resultid="2291" swimtime="00:03:53.55"><SPLITS><SPLIT distance="50" swimtime="00:00:49.22"/><SPLIT distance="100" swimtime="00:01:47.94"/><SPLIT distance="150" swimtime="00:02:49.95"/></SPLITS></RESULT><RESULT eventid="32" heatid="346" lane="2" points="116" resultid="2576" swimtime="00:01:56.44"><SPLITS><SPLIT distance="50" swimtime="00:00:55.06"/></SPLITS></RESULT><RESULT eventid="40" heatid="453" lane="2" resultid="3383" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="208" birthdate="2015-01-01" firstname="Samuel" gender="M" lastname="Weber" license="482343"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="28" lane="4" points="88" resultid="208" swimtime="00:00:58.29"><SPLITS/></RESULT><RESULT eventid="10" heatid="135" lane="2" points="77" resultid="1014" swimtime="00:00:49.06"><SPLITS/></RESULT><RESULT eventid="14" heatid="210" lane="1" points="72" resultid="1590" swimtime="00:02:04.01"><SPLITS><SPLIT distance="50" swimtime="00:01:00.62"/></SPLITS></RESULT><RESULT eventid="28" heatid="276" lane="4" points="77" resultid="2050" swimtime="00:00:55.66"><SPLITS/></RESULT><RESULT eventid="32" heatid="346" lane="7" points="82" resultid="2580" swimtime="00:02:10.45"><SPLITS><SPLIT distance="50" swimtime="00:00:59.35"/></SPLITS></RESULT><RESULT eventid="40" heatid="452" lane="2" points="67" resultid="3375" swimtime="00:01:55.06"><SPLITS><SPLIT distance="50" swimtime="00:00:52.12"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="212" birthdate="2014-01-01" firstname="Lucas" gender="M" lastname="Song" license="449255"><HANDICAP/><ENTRIES/><RESULTS><RESULT comment="09:41 Start vor dem Startsignal" eventid="2" heatid="28" lane="8" resultid="212" status="DSQ" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="10" heatid="136" lane="5" points="102" resultid="1025" swimtime="00:00:44.67"><SPLITS/></RESULT><RESULT eventid="14" heatid="213" lane="3" points="98" resultid="1615" swimtime="00:01:51.86"><SPLITS><SPLIT distance="50" swimtime="00:00:55.57"/></SPLITS></RESULT><RESULT eventid="28" heatid="277" lane="3" points="104" resultid="2056" swimtime="00:00:50.30"><SPLITS/></RESULT><RESULT eventid="40" heatid="453" lane="6" points="96" resultid="3387" swimtime="00:01:42.15"><SPLITS><SPLIT distance="50" swimtime="00:00:46.12"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="214" birthdate="2014-01-01" firstname="Florian" gender="M" lastname="Aign" license="449247"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="29" lane="2" points="136" resultid="214" swimtime="00:00:50.39"><SPLITS/></RESULT><RESULT eventid="8" heatid="93" lane="2" points="139" resultid="698" swimtime="00:04:03.10"><SPLITS><SPLIT distance="50" swimtime="00:00:53.74"/><SPLIT distance="100" swimtime="00:01:56.06"/><SPLIT distance="150" swimtime="00:03:01.06"/></SPLITS></RESULT><RESULT eventid="10" heatid="138" lane="8" points="162" resultid="1043" swimtime="00:00:38.34"><SPLITS/></RESULT><RESULT eventid="14" heatid="215" lane="2" points="124" resultid="1629" swimtime="00:01:43.21"><SPLITS><SPLIT distance="50" swimtime="00:00:52.65"/></SPLITS></RESULT><RESULT eventid="30" heatid="311" lane="3" points="141" resultid="2314" swimtime="00:03:15.60"><SPLITS><SPLIT distance="50" swimtime="00:00:41.77"/><SPLIT distance="100" swimtime="00:01:31.46"/><SPLIT distance="150" swimtime="00:02:26.46"/></SPLITS></RESULT><RESULT eventid="32" heatid="348" lane="7" points="132" resultid="2596" swimtime="00:01:51.64"><SPLITS><SPLIT distance="50" swimtime="00:00:53.30"/></SPLITS></RESULT><RESULT eventid="38" heatid="414" lane="2" points="135" resultid="3084" swimtime="00:03:38.09"><SPLITS><SPLIT distance="50" swimtime="00:00:52.49"/><SPLIT distance="100" swimtime="00:01:47.74"/><SPLIT distance="150" swimtime="00:02:44.71"/></SPLITS></RESULT><RESULT eventid="40" heatid="457" lane="1" points="137" resultid="3413" swimtime="00:01:30.76"><SPLITS><SPLIT distance="50" swimtime="00:00:42.35"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="218" birthdate="2013-01-01" firstname="Darwin" gender="M" lastname="Koch" license="443857"><HANDICAP/><ENTRIES/><RESULTS><RESULT comment="09:42 Start vor dem Startsignal" eventid="2" heatid="29" lane="6" resultid="218" status="DSQ" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="8" heatid="94" lane="1" points="156" resultid="704" swimtime="00:03:53.67"><SPLITS><SPLIT distance="50" swimtime="00:00:56.29"/><SPLIT distance="100" swimtime="00:01:55.24"/><SPLIT distance="150" swimtime="00:02:56.70"/></SPLITS></RESULT><RESULT eventid="10" heatid="137" lane="5" points="136" resultid="1033" swimtime="00:00:40.66"><SPLITS/></RESULT><RESULT eventid="14" heatid="213" lane="1" points="130" resultid="1613" swimtime="00:01:41.70"><SPLITS><SPLIT distance="50" swimtime="00:00:49.98"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="244" birthdate="2014-01-01" firstname="Arvin Mateo" gender="M" lastname="Azadeh Reimondez" license="449261"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="32" lane="8" points="129" resultid="244" swimtime="00:00:51.34"><SPLITS/></RESULT><RESULT eventid="8" heatid="94" lane="6" points="145" resultid="709" swimtime="00:03:59.52"><SPLITS><SPLIT distance="50" swimtime="00:00:55.13"/><SPLIT distance="100" swimtime="00:01:57.27"/><SPLIT distance="150" swimtime="00:03:01.06"/></SPLITS></RESULT><RESULT eventid="10" heatid="137" lane="7" points="112" resultid="1035" swimtime="00:00:43.27"><SPLITS/></RESULT><RESULT eventid="14" heatid="211" lane="1" points="92" resultid="1598" swimtime="00:01:54.15"><SPLITS><SPLIT distance="50" swimtime="00:00:58.11"/></SPLITS></RESULT><RESULT eventid="28" heatid="275" lane="3" points="107" resultid="2041" swimtime="00:00:49.88"><SPLITS/></RESULT><RESULT eventid="30" heatid="309" lane="4" points="94" resultid="2299" swimtime="00:03:43.97"><SPLITS><SPLIT distance="50" swimtime="00:00:51.16"/><SPLIT distance="100" swimtime="00:01:50.38"/><SPLIT distance="150" swimtime="00:02:48.90"/></SPLITS></RESULT><RESULT eventid="32" heatid="347" lane="5" points="113" resultid="2586" swimtime="00:01:57.61"><SPLITS><SPLIT distance="50" swimtime="00:00:57.54"/></SPLITS></RESULT><RESULT eventid="40" heatid="454" lane="5" points="98" resultid="3394" swimtime="00:01:41.56"><SPLITS><SPLIT distance="50" swimtime="00:00:49.31"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="246" birthdate="2013-01-01" firstname="Kilian" gender="M" lastname="Sußbauer" license="445749"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="33" lane="2" points="179" resultid="246" swimtime="00:00:45.97"><SPLITS/></RESULT><RESULT eventid="8" heatid="97" lane="6" points="223" resultid="731" swimtime="00:03:27.48"><SPLITS><SPLIT distance="50" swimtime="00:00:49.30"/><SPLIT distance="100" swimtime="00:01:42.15"/><SPLIT distance="150" swimtime="00:02:37.04"/></SPLITS></RESULT><RESULT eventid="10" heatid="140" lane="4" points="176" resultid="1055" swimtime="00:00:37.31"><SPLITS/></RESULT><RESULT eventid="12" heatid="179" lane="5" points="213" resultid="1354" swimtime="00:03:10.61"><SPLITS><SPLIT distance="50" swimtime="00:00:47.74"/><SPLIT distance="100" swimtime="00:01:35.79"/><SPLIT distance="150" swimtime="00:02:27.90"/></SPLITS></RESULT><RESULT eventid="30" heatid="314" lane="4" points="194" resultid="2337" swimtime="00:02:56.02"><SPLITS><SPLIT distance="50" swimtime="00:00:40.64"/><SPLIT distance="100" swimtime="00:01:27.43"/><SPLIT distance="150" swimtime="00:02:13.86"/></SPLITS></RESULT><RESULT eventid="32" heatid="350" lane="3" points="197" resultid="2607" swimtime="00:01:37.74"><SPLITS><SPLIT distance="50" swimtime="00:00:46.88"/></SPLITS></RESULT><RESULT eventid="36" heatid="387" lane="4" points="122" resultid="2881" swimtime="00:00:44.83"><SPLITS/></RESULT><RESULT eventid="40" heatid="460" lane="3" points="183" resultid="3438" swimtime="00:01:22.46"><SPLITS><SPLIT distance="50" swimtime="00:00:39.99"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="250" birthdate="2013-01-01" firstname="Maximilian" gender="M" lastname="Meier" license="462715"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="33" lane="6" points="215" resultid="250" swimtime="00:00:43.29"><SPLITS/></RESULT><RESULT eventid="8" heatid="97" lane="3" points="244" resultid="728" swimtime="00:03:21.50"><SPLITS><SPLIT distance="50" swimtime="00:00:46.46"/><SPLIT distance="100" swimtime="00:01:40.02"/><SPLIT distance="150" swimtime="00:02:32.57"/></SPLITS></RESULT><RESULT eventid="10" heatid="141" lane="4" points="227" resultid="1062" swimtime="00:00:34.24"><SPLITS/></RESULT><RESULT eventid="14" heatid="212" lane="7" points="221" resultid="1611" swimtime="00:01:25.31"><SPLITS><SPLIT distance="50" swimtime="00:00:41.44"/></SPLITS></RESULT><RESULT eventid="28" heatid="279" lane="7" points="207" resultid="2075" swimtime="00:00:40.05"><SPLITS/></RESULT><RESULT eventid="30" heatid="315" lane="2" points="241" resultid="2343" swimtime="00:02:43.78"><SPLITS><SPLIT distance="50" swimtime="00:00:37.10"/><SPLIT distance="100" swimtime="00:01:19.75"/><SPLIT distance="150" swimtime="00:02:03.35"/></SPLITS></RESULT><RESULT eventid="36" heatid="385" lane="2" points="142" resultid="2864" swimtime="00:00:42.68"><SPLITS/></RESULT><RESULT eventid="40" heatid="463" lane="8" points="232" resultid="3466" swimtime="00:01:16.16"><SPLITS><SPLIT distance="50" swimtime="00:00:36.94"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="269" birthdate="2013-01-01" firstname="Paul" gender="M" lastname="Nowey" license="443841"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="36" lane="3" points="257" resultid="269" swimtime="00:00:40.80"><SPLITS/></RESULT><RESULT eventid="8" heatid="99" lane="6" points="349" resultid="746" swimtime="00:02:58.85"><SPLITS><SPLIT distance="50" swimtime="00:00:40.77"/><SPLIT distance="100" swimtime="00:01:26.84"/><SPLIT distance="150" swimtime="00:02:12.94"/></SPLITS></RESULT><RESULT eventid="10" heatid="144" lane="8" points="236" resultid="1089" swimtime="00:00:33.83"><SPLITS/></RESULT><RESULT eventid="12" heatid="183" lane="6" points="295" resultid="1387" swimtime="00:02:51.09"><SPLITS><SPLIT distance="50" swimtime="00:00:38.55"/><SPLIT distance="100" swimtime="00:01:26.91"/><SPLIT distance="150" swimtime="00:02:11.98"/></SPLITS></RESULT><RESULT eventid="26" heatid="251" lane="2" resultid="1856" swimtime="00:00:53.16"><SPLITS/></RESULT><RESULT eventid="30" heatid="318" lane="2" points="247" resultid="2367" swimtime="00:02:42.41"><SPLITS><SPLIT distance="50" swimtime="00:00:37.33"/><SPLIT distance="100" swimtime="00:01:19.11"/><SPLIT distance="150" swimtime="00:02:02.16"/></SPLITS></RESULT><RESULT eventid="32" heatid="353" lane="8" points="290" resultid="2634" swimtime="00:01:25.92"><SPLITS><SPLIT distance="50" swimtime="00:00:41.29"/></SPLITS></RESULT><RESULT eventid="38" heatid="413" lane="7" points="217" resultid="3082" swimtime="00:03:06.10"><SPLITS><SPLIT distance="50" swimtime="00:00:42.80"/><SPLIT distance="100" swimtime="00:01:31.58"/><SPLIT distance="150" swimtime="00:02:19.09"/></SPLITS></RESULT><RESULT eventid="40" heatid="464" lane="5" points="248" resultid="3471" swimtime="00:01:14.50"><SPLITS><SPLIT distance="50" swimtime="00:00:35.74"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="271" birthdate="2011-01-01" firstname="Franz" gender="M" lastname="Rummel" license="431792"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="36" lane="5" points="287" resultid="271" swimtime="00:00:39.32"><SPLITS/></RESULT><RESULT eventid="10" heatid="147" lane="5" points="321" resultid="1110" swimtime="00:00:30.51"><SPLITS/></RESULT><RESULT eventid="12" heatid="185" lane="6" points="337" resultid="1401" swimtime="00:02:43.81"><SPLITS><SPLIT distance="50" swimtime="00:00:35.26"/><SPLIT distance="100" swimtime="00:01:18.95"/><SPLIT distance="150" swimtime="00:02:06.62"/></SPLITS></RESULT><RESULT eventid="30" heatid="320" lane="6" points="361" resultid="2387" swimtime="00:02:23.24"><SPLITS><SPLIT distance="50" swimtime="00:00:31.86"/><SPLIT distance="100" swimtime="00:01:08.37"/><SPLIT distance="150" swimtime="00:01:46.45"/></SPLITS></RESULT><RESULT eventid="32" heatid="352" lane="5" points="258" resultid="2623" swimtime="00:01:29.27"><SPLITS><SPLIT distance="50" swimtime="00:00:41.17"/></SPLITS></RESULT><RESULT eventid="36" heatid="392" lane="4" points="283" resultid="2921" swimtime="00:00:33.90"><SPLITS/></RESULT><RESULT eventid="40" heatid="467" lane="4" points="333" resultid="3493" swimtime="00:01:07.55"><SPLITS><SPLIT distance="50" swimtime="00:00:31.91"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="302" birthdate="2009-01-01" firstname="Dimitar" gender="M" lastname="Todorovski" license="478501"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="40" lane="4" points="549" resultid="302" swimtime="00:00:31.68"><SPLITS/></RESULT><RESULT eventid="8" heatid="101" lane="3" points="511" resultid="759" swimtime="00:02:37.49"><SPLITS><SPLIT distance="50" swimtime="00:00:35.26"/><SPLIT distance="100" swimtime="00:01:15.88"/><SPLIT distance="150" swimtime="00:01:57.42"/></SPLITS></RESULT><RESULT eventid="10" heatid="153" lane="4" points="431" resultid="1157" swimtime="00:00:27.67"><SPLITS/></RESULT><RESULT eventid="32" heatid="356" lane="5" points="495" resultid="2654" swimtime="00:01:11.89"><SPLITS><SPLIT distance="50" swimtime="00:00:33.18"/></SPLITS></RESULT><RESULT eventid="36" heatid="396" lane="3" points="426" resultid="2952" swimtime="00:00:29.59"><SPLITS/></RESULT><RESULT eventid="40" heatid="472" lane="7" points="487" resultid="3536" swimtime="00:00:59.53"><SPLITS><SPLIT distance="50" swimtime="00:00:27.77"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="304" birthdate="2009-01-01" firstname="Damjan" gender="M" lastname="Todorovski" license="478502"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="40" lane="6" points="505" resultid="304" swimtime="00:00:32.58"><SPLITS/></RESULT><RESULT eventid="8" heatid="101" lane="7" points="449" resultid="762" swimtime="00:02:44.46"><SPLITS><SPLIT distance="50" swimtime="00:00:34.95"/><SPLIT distance="100" swimtime="00:01:18.14"/><SPLIT distance="150" swimtime="00:02:01.49"/></SPLITS></RESULT><RESULT eventid="10" heatid="151" lane="3" points="344" resultid="1140" swimtime="00:00:29.84"><SPLITS/></RESULT><RESULT eventid="32" heatid="356" lane="2" points="466" resultid="2651" swimtime="00:01:13.34"><SPLITS><SPLIT distance="50" swimtime="00:00:33.05"/></SPLITS></RESULT><RESULT eventid="36" heatid="396" lane="2" points="406" resultid="2951" swimtime="00:00:30.07"><SPLITS/></RESULT><RESULT eventid="40" heatid="471" lane="8" points="402" resultid="3529" swimtime="00:01:03.49"><SPLITS><SPLIT distance="50" swimtime="00:00:30.29"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="339" birthdate="2014-01-01" firstname="Jovana" gender="F" lastname="Todorovska" license="478503"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="46" lane="7" points="298" resultid="350" swimtime="00:05:53.59"><SPLITS><SPLIT distance="100" swimtime="00:01:22.66"/><SPLIT distance="200" swimtime="00:02:53.66"/><SPLIT distance="300" swimtime="00:04:26.31"/></SPLITS></RESULT><RESULT eventid="11" heatid="169" lane="8" points="341" resultid="1282" swimtime="00:03:00.51"><SPLITS><SPLIT distance="50" swimtime="00:00:40.64"/><SPLIT distance="100" swimtime="00:01:26.04"/><SPLIT distance="150" swimtime="00:02:20.77"/></SPLITS></RESULT><RESULT eventid="13" heatid="204" lane="7" points="301" resultid="1550" swimtime="00:01:25.71"><SPLITS><SPLIT distance="50" swimtime="00:00:41.67"/></SPLITS></RESULT><RESULT eventid="19" heatid="235" lane="3" resultid="1764" swimtime="00:00:53.99"><SPLITS/></RESULT><RESULT eventid="21" heatid="238" lane="3" resultid="1780" swimtime="00:00:53.52"><SPLITS/></RESULT><RESULT eventid="29" heatid="299" lane="8" points="284" resultid="2229" swimtime="00:02:51.87"><SPLITS><SPLIT distance="50" swimtime="00:00:38.18"/><SPLIT distance="100" swimtime="00:01:22.87"/><SPLIT distance="150" swimtime="00:02:08.64"/></SPLITS></RESULT><RESULT eventid="37" heatid="407" lane="4" points="321" resultid="3034" swimtime="00:03:00.13"><SPLITS><SPLIT distance="50" swimtime="00:00:41.60"/><SPLIT distance="100" swimtime="00:01:28.15"/><SPLIT distance="150" swimtime="00:02:15.13"/></SPLITS></RESULT><RESULT eventid="39" heatid="438" lane="2" points="343" resultid="3267" swimtime="00:01:13.87"><SPLITS><SPLIT distance="50" swimtime="00:00:35.20"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="345" birthdate="2012-01-01" firstname="Helene" gender="F" lastname="Herdeg" license="443834"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="48" lane="4" points="391" resultid="362" swimtime="00:05:23.20"><SPLITS><SPLIT distance="100" swimtime="00:01:17.57"/><SPLIT distance="200" swimtime="00:02:42.12"/><SPLIT distance="300" swimtime="00:04:06.00"/></SPLITS></RESULT><RESULT eventid="9" heatid="119" lane="5" points="361" resultid="900" swimtime="00:00:33.24"><SPLITS/></RESULT><RESULT eventid="11" heatid="168" lane="8" points="341" resultid="1274" swimtime="00:03:00.52"><SPLITS><SPLIT distance="50" swimtime="00:00:41.63"/><SPLIT distance="100" swimtime="00:01:27.99"/><SPLIT distance="150" swimtime="00:02:21.75"/></SPLITS></RESULT><RESULT eventid="29" heatid="301" lane="4" points="403" resultid="2240" swimtime="00:02:32.94"><SPLITS><SPLIT distance="50" swimtime="00:00:34.48"/><SPLIT distance="100" swimtime="00:01:14.24"/><SPLIT distance="150" swimtime="00:01:54.70"/></SPLITS></RESULT><RESULT eventid="35" heatid="368" lane="2" points="264" resultid="2736" swimtime="00:00:38.08"><SPLITS/></RESULT><RESULT eventid="39" heatid="439" lane="4" points="384" resultid="3277" swimtime="00:01:11.13"><SPLITS><SPLIT distance="50" swimtime="00:00:33.77"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="352" birthdate="2011-01-01" firstname="Lina" gender="F" lastname="Sinkel" license="424441"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="49" lane="3" points="394" resultid="369" swimtime="00:05:22.44"><SPLITS><SPLIT distance="100" swimtime="00:01:15.05"/><SPLIT distance="200" swimtime="00:02:38.41"/><SPLIT distance="300" swimtime="00:04:02.26"/></SPLITS></RESULT><RESULT eventid="9" heatid="122" lane="6" points="420" resultid="925" swimtime="00:00:31.60"><SPLITS/></RESULT><RESULT eventid="13" heatid="204" lane="3" points="360" resultid="1546" swimtime="00:01:20.75"><SPLITS><SPLIT distance="50" swimtime="00:00:38.56"/></SPLITS></RESULT><RESULT eventid="29" heatid="303" lane="6" points="431" resultid="2258" swimtime="00:02:29.52"><SPLITS><SPLIT distance="50" swimtime="00:00:34.03"/><SPLIT distance="100" swimtime="00:01:12.58"/><SPLIT distance="150" swimtime="00:01:50.84"/></SPLITS></RESULT><RESULT eventid="35" heatid="375" lane="4" points="379" resultid="2793" swimtime="00:00:33.73"><SPLITS/></RESULT><RESULT eventid="37" heatid="407" lane="5" points="356" resultid="3035" swimtime="00:02:53.95"><SPLITS><SPLIT distance="50" swimtime="00:00:40.58"/><SPLIT distance="100" swimtime="00:01:24.50"/><SPLIT distance="150" swimtime="00:02:09.36"/></SPLITS></RESULT><RESULT eventid="39" heatid="442" lane="8" points="417" resultid="3304" swimtime="00:01:09.20"><SPLITS><SPLIT distance="50" swimtime="00:00:33.52"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="364" birthdate="2010-01-01" firstname="Mia" gender="F" lastname="Mahl" license="414341"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="51" lane="1" points="450" resultid="383" swimtime="00:05:08.33"><SPLITS><SPLIT distance="100" swimtime="00:01:11.74"/><SPLIT distance="200" swimtime="00:02:31.93"/><SPLIT distance="300" swimtime="00:03:51.31"/></SPLITS></RESULT><RESULT eventid="9" heatid="125" lane="4" points="472" resultid="947" swimtime="00:00:30.38"><SPLITS/></RESULT><RESULT eventid="11" heatid="171" lane="2" points="456" resultid="1292" swimtime="00:02:43.75"><SPLITS><SPLIT distance="50" swimtime="00:00:35.75"/><SPLIT distance="100" swimtime="00:01:16.47"/><SPLIT distance="150" swimtime="00:02:07.18"/></SPLITS></RESULT><RESULT eventid="13" heatid="205" lane="3" points="415" resultid="1554" swimtime="00:01:16.96"><SPLITS><SPLIT distance="50" swimtime="00:00:37.37"/></SPLITS></RESULT><RESULT eventid="27" heatid="268" lane="6" points="424" resultid="1993" swimtime="00:00:35.90"><SPLITS/></RESULT><RESULT eventid="29" heatid="305" lane="7" points="487" resultid="2273" swimtime="00:02:23.52"><SPLITS><SPLIT distance="50" swimtime="00:00:32.22"/><SPLIT distance="100" swimtime="00:01:08.57"/><SPLIT distance="150" swimtime="00:01:45.85"/></SPLITS></RESULT><RESULT eventid="37" heatid="409" lane="4" points="415" resultid="3050" swimtime="00:02:45.30"><SPLITS><SPLIT distance="50" swimtime="00:00:37.65"/><SPLIT distance="100" swimtime="00:01:20.10"/><SPLIT distance="150" swimtime="00:02:03.66"/></SPLITS></RESULT><RESULT eventid="39" heatid="447" lane="8" points="472" resultid="3342" swimtime="00:01:06.39"><SPLITS><SPLIT distance="50" swimtime="00:00:32.16"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="366" birthdate="2012-01-01" firstname="Emma" gender="F" lastname="Irrgang" license="443835"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="51" lane="4" points="496" resultid="385" swimtime="00:04:58.50"><SPLITS><SPLIT distance="100" swimtime="00:01:09.00"/><SPLIT distance="200" swimtime="00:02:27.76"/></SPLITS></RESULT><RESULT eventid="5" heatid="70" lane="8" points="438" resultid="527" swimtime="00:01:13.01"><SPLITS><SPLIT distance="50" swimtime="00:00:33.96"/></SPLITS></RESULT><RESULT eventid="11" heatid="173" lane="1" points="496" resultid="1307" swimtime="00:02:39.30"><SPLITS><SPLIT distance="50" swimtime="00:00:34.32"/><SPLIT distance="100" swimtime="00:01:16.46"/><SPLIT distance="150" swimtime="00:02:03.97"/></SPLITS></RESULT><RESULT eventid="29" heatid="306" lane="8" points="547" resultid="2282" swimtime="00:02:18.07"><SPLITS><SPLIT distance="50" swimtime="00:00:32.98"/><SPLIT distance="100" swimtime="00:01:08.84"/><SPLIT distance="150" swimtime="00:01:44.31"/></SPLITS></RESULT><RESULT eventid="35" heatid="379" lane="6" points="424" resultid="2825" swimtime="00:00:32.51"><SPLITS/></RESULT><RESULT eventid="39" heatid="448" lane="6" points="531" resultid="3348" swimtime="00:01:03.85"><SPLITS><SPLIT distance="50" swimtime="00:00:30.65"/></SPLITS></RESULT><RESULT eventid="41" heatid="477" lane="5" points="474" resultid="3567" swimtime="00:05:41.43"><SPLITS><SPLIT distance="50" swimtime="00:00:35.67"/><SPLIT distance="100" swimtime="00:01:19.00"/><SPLIT distance="150" swimtime="00:02:01.87"/><SPLIT distance="200" swimtime="00:02:43.59"/><SPLIT distance="250" swimtime="00:03:32.83"/><SPLIT distance="300" swimtime="00:04:24.82"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="370" birthdate="2006-01-01" firstname="Amira" gender="F" lastname="Varna" license="358238"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="51" lane="8" points="452" resultid="389" swimtime="00:05:07.84"><SPLITS><SPLIT distance="100" swimtime="00:01:11.03"/><SPLIT distance="200" swimtime="00:02:29.67"/><SPLIT distance="300" swimtime="00:03:49.34"/></SPLITS></RESULT><RESULT eventid="9" heatid="129" lane="2" points="495" resultid="976" swimtime="00:00:29.92"><SPLITS/></RESULT><RESULT eventid="29" heatid="305" lane="6" points="509" resultid="2272" swimtime="00:02:21.43"><SPLITS><SPLIT distance="50" swimtime="00:00:32.31"/><SPLIT distance="100" swimtime="00:01:07.83"/><SPLIT distance="150" swimtime="00:01:44.98"/></SPLITS></RESULT><RESULT eventid="39" heatid="448" lane="7" points="517" resultid="3349" swimtime="00:01:04.39"><SPLITS><SPLIT distance="50" swimtime="00:00:30.91"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="401" birthdate="2014-01-01" firstname="Michael" gender="M" lastname="Ustyuzhaninov" license="449266"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="57" lane="2" points="241" resultid="427" swimtime="00:05:53.44"><SPLITS><SPLIT distance="100" swimtime="00:01:21.15"/><SPLIT distance="200" swimtime="00:02:53.47"/><SPLIT distance="300" swimtime="00:04:24.87"/></SPLITS></RESULT><RESULT eventid="8" heatid="98" lane="1" points="269" resultid="734" swimtime="00:03:14.96"><SPLITS><SPLIT distance="50" swimtime="00:00:45.40"/><SPLIT distance="100" swimtime="00:01:34.42"/><SPLIT distance="150" swimtime="00:02:26.67"/></SPLITS></RESULT><RESULT eventid="12" heatid="179" lane="1" points="234" resultid="1350" swimtime="00:03:04.99"><SPLITS><SPLIT distance="50" swimtime="00:00:40.74"/><SPLIT distance="100" swimtime="00:01:33.27"/><SPLIT distance="150" swimtime="00:02:24.49"/></SPLITS></RESULT><RESULT eventid="26" heatid="251" lane="3" resultid="1857" swimtime="00:00:54.23"><SPLITS/></RESULT><RESULT eventid="32" heatid="351" lane="1" points="238" resultid="2612" swimtime="00:01:31.76"><SPLITS><SPLIT distance="50" swimtime="00:00:43.87"/></SPLITS></RESULT><RESULT eventid="36" heatid="388" lane="8" points="155" resultid="2893" swimtime="00:00:41.43"><SPLITS/></RESULT><RESULT eventid="40" heatid="462" lane="1" points="201" resultid="3452" swimtime="00:01:19.95"><SPLITS><SPLIT distance="50" swimtime="00:00:38.16"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="417" birthdate="2012-01-01" firstname="Maxim" gender="M" lastname="Belyaev" license="442808"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="59" lane="6" points="299" resultid="446" swimtime="00:05:28.99"><SPLITS><SPLIT distance="100" swimtime="00:01:16.24"/><SPLIT distance="200" swimtime="00:02:40.31"/><SPLIT distance="300" swimtime="00:04:06.06"/></SPLITS></RESULT><RESULT eventid="10" heatid="147" lane="7" points="297" resultid="1112" swimtime="00:00:31.32"><SPLITS/></RESULT><RESULT eventid="12" heatid="184" lane="3" points="313" resultid="1391" swimtime="00:02:47.80"><SPLITS><SPLIT distance="50" swimtime="00:00:36.29"/><SPLIT distance="100" swimtime="00:01:19.61"/><SPLIT distance="150" swimtime="00:02:10.81"/></SPLITS></RESULT><RESULT eventid="14" heatid="222" lane="8" points="309" resultid="1689" swimtime="00:01:16.25"><SPLITS><SPLIT distance="50" swimtime="00:00:37.30"/></SPLITS></RESULT><RESULT eventid="30" heatid="320" lane="5" points="326" resultid="2386" swimtime="00:02:28.19"><SPLITS><SPLIT distance="50" swimtime="00:01:50.71"/><SPLIT distance="100" swimtime="00:01:10.96"/></SPLITS></RESULT><RESULT eventid="38" heatid="417" lane="5" points="313" resultid="3111" swimtime="00:02:44.81"><SPLITS><SPLIT distance="50" swimtime="00:00:37.56"/><SPLIT distance="100" swimtime="00:01:19.65"/><SPLIT distance="150" swimtime="00:02:02.33"/></SPLITS></RESULT><RESULT eventid="40" heatid="466" lane="4" points="281" resultid="3486" swimtime="00:01:11.51"><SPLITS><SPLIT distance="50" swimtime="00:00:33.51"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="421" birthdate="2011-01-01" firstname="Marc" gender="M" lastname="Rohrmüller" license="424439"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="60" lane="2" points="401" resultid="450" swimtime="00:04:58.25"><SPLITS><SPLIT distance="100" swimtime="00:01:11.29"/><SPLIT distance="200" swimtime="00:02:27.55"/><SPLIT distance="300" swimtime="00:03:46.18"/></SPLITS></RESULT><RESULT eventid="10" heatid="150" lane="6" points="403" resultid="1135" swimtime="00:00:28.29"><SPLITS/></RESULT><RESULT eventid="36" heatid="395" lane="1" points="371" resultid="2942" swimtime="00:00:30.98"><SPLITS/></RESULT><RESULT eventid="40" heatid="469" lane="5" points="458" resultid="3510" swimtime="00:01:00.76"><SPLITS><SPLIT distance="50" swimtime="00:00:29.81"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="425" birthdate="2011-01-01" firstname="Raúl" gender="M" lastname="Muñoz" license="424436"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="60" lane="7" points="401" resultid="454" swimtime="00:04:58.25"><SPLITS><SPLIT distance="100" swimtime="00:01:09.78"/><SPLIT distance="200" swimtime="00:02:26.53"/><SPLIT distance="300" swimtime="00:03:45.39"/></SPLITS></RESULT><RESULT eventid="10" heatid="148" lane="6" points="353" resultid="1119" swimtime="00:00:29.56"><SPLITS/></RESULT><RESULT eventid="14" heatid="222" lane="2" points="269" resultid="1683" swimtime="00:01:19.85"><SPLITS><SPLIT distance="50" swimtime="00:00:38.65"/></SPLITS></RESULT><RESULT eventid="30" heatid="322" lane="1" points="392" resultid="2396" swimtime="00:02:19.26"><SPLITS><SPLIT distance="50" swimtime="00:00:32.25"/><SPLIT distance="100" swimtime="00:01:07.75"/><SPLIT distance="150" swimtime="00:01:44.66"/></SPLITS></RESULT><RESULT eventid="36" heatid="392" lane="7" points="202" resultid="2924" swimtime="00:00:37.94"><SPLITS/></RESULT><RESULT eventid="40" heatid="468" lane="4" points="380" resultid="3501" swimtime="00:01:04.64"><SPLITS><SPLIT distance="50" swimtime="00:00:31.47"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="429" birthdate="2010-01-01" firstname="Andrew" gender="M" lastname="Cicero" license="412140"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="61" lane="3" points="484" resultid="458" swimtime="00:04:40.12"><SPLITS><SPLIT distance="100" swimtime="00:01:03.72"/><SPLIT distance="200" swimtime="00:02:15.15"/><SPLIT distance="300" swimtime="00:03:28.47"/></SPLITS></RESULT><RESULT eventid="12" heatid="187" lane="3" points="419" resultid="1414" swimtime="00:02:32.30"><SPLITS><SPLIT distance="50" swimtime="00:00:33.36"/><SPLIT distance="100" swimtime="00:01:09.85"/><SPLIT distance="150" swimtime="00:02:00.14"/></SPLITS></RESULT><RESULT eventid="18" heatid="232" lane="5" points="475" resultid="1751" swimtime="00:09:39.19"><SPLITS><SPLIT distance="100" swimtime="00:01:06.21"/><SPLIT distance="200" swimtime="00:02:18.71"/><SPLIT distance="300" swimtime="00:03:31.61"/><SPLIT distance="400" swimtime="00:04:45.14"/><SPLIT distance="500" swimtime="00:05:59.26"/><SPLIT distance="600" swimtime="00:07:14.06"/><SPLIT distance="700" swimtime="00:08:28.18"/></SPLITS></RESULT><RESULT eventid="30" heatid="323" lane="2" points="459" resultid="2405" swimtime="00:02:12.17"><SPLITS><SPLIT distance="50" swimtime="00:00:30.07"/><SPLIT distance="100" swimtime="00:01:04.40"/><SPLIT distance="150" swimtime="00:01:38.41"/></SPLITS></RESULT><RESULT eventid="38" heatid="419" lane="1" points="429" resultid="3121" swimtime="00:02:28.37"><SPLITS><SPLIT distance="50" swimtime="00:00:34.92"/><SPLIT distance="100" swimtime="00:01:13.43"/><SPLIT distance="150" swimtime="00:01:52.31"/></SPLITS></RESULT><RESULT eventid="42" heatid="480" lane="1" points="423" resultid="3585" swimtime="00:05:24.62"><SPLITS><SPLIT distance="50" swimtime="00:00:35.56"/><SPLIT distance="100" swimtime="00:01:18.57"/><SPLIT distance="150" swimtime="00:01:57.77"/><SPLIT distance="200" swimtime="00:02:36.90"/><SPLIT distance="250" swimtime="00:03:28.79"/><SPLIT distance="300" swimtime="00:04:18.24"/><SPLIT distance="350" swimtime="00:04:51.95"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="441" birthdate="2013-01-01" firstname="Linda" gender="F" lastname="Mahl" license="443844"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="5" heatid="64" lane="4" points="196" resultid="476" swimtime="00:01:35.49"><SPLITS><SPLIT distance="50" swimtime="00:00:41.39"/></SPLITS></RESULT><RESULT eventid="7" heatid="88" lane="4" points="331" resultid="660" swimtime="00:03:20.69"><SPLITS><SPLIT distance="50" swimtime="00:00:46.53"/><SPLIT distance="100" swimtime="00:01:39.33"/><SPLIT distance="150" swimtime="00:02:29.64"/></SPLITS></RESULT><RESULT eventid="9" heatid="115" lane="2" points="305" resultid="866" swimtime="00:00:35.13"><SPLITS/></RESULT><RESULT eventid="13" heatid="198" lane="3" points="252" resultid="1498" swimtime="00:01:30.95"><SPLITS><SPLIT distance="50" swimtime="00:00:44.88"/></SPLITS></RESULT><RESULT eventid="21" heatid="238" lane="2" resultid="1779" swimtime="00:00:59.14"><SPLITS/></RESULT><RESULT eventid="29" heatid="298" lane="2" points="310" resultid="2215" swimtime="00:02:46.86"><SPLITS><SPLIT distance="50" swimtime="00:00:38.42"/><SPLIT distance="100" swimtime="00:01:20.43"/><SPLIT distance="150" swimtime="00:02:04.87"/></SPLITS></RESULT><RESULT eventid="31" heatid="339" lane="2" points="355" resultid="2524" swimtime="00:01:30.52"><SPLITS><SPLIT distance="50" swimtime="00:00:42.65"/></SPLITS></RESULT><RESULT eventid="35" heatid="369" lane="5" points="218" resultid="2747" swimtime="00:00:40.53"><SPLITS/></RESULT><RESULT eventid="39" heatid="435" lane="1" points="308" resultid="3242" swimtime="00:01:16.49"><SPLITS><SPLIT distance="50" swimtime="00:00:37.58"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="452" birthdate="2013-01-01" firstname="Valentina" gender="F" lastname="Rößger" license="443851"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="5" heatid="67" lane="7" points="267" resultid="502" swimtime="00:01:26.10"><SPLITS><SPLIT distance="50" swimtime="00:00:36.70"/></SPLITS></RESULT><RESULT eventid="7" heatid="88" lane="1" points="329" resultid="657" swimtime="00:03:21.14"><SPLITS><SPLIT distance="50" swimtime="00:00:46.55"/><SPLIT distance="100" swimtime="00:01:37.14"/><SPLIT distance="150" swimtime="00:02:30.65"/></SPLITS></RESULT><RESULT eventid="9" heatid="125" lane="3" points="466" resultid="946" swimtime="00:00:30.53"><SPLITS/></RESULT><RESULT eventid="11" heatid="169" lane="2" points="384" resultid="1276" swimtime="00:02:53.44"><SPLITS><SPLIT distance="50" swimtime="00:00:37.07"/><SPLIT distance="100" swimtime="00:01:23.22"/><SPLIT distance="150" swimtime="00:02:15.57"/></SPLITS></RESULT><RESULT eventid="21" heatid="238" lane="5" resultid="1782" swimtime="00:00:47.24"><SPLITS/></RESULT><RESULT eventid="23" heatid="243" lane="5" resultid="1811" swimtime="00:00:50.71"><SPLITS/></RESULT><RESULT eventid="29" heatid="300" lane="4" points="359" resultid="2233" swimtime="00:02:38.83"><SPLITS><SPLIT distance="50" swimtime="00:00:34.81"/><SPLIT distance="100" swimtime="00:01:15.93"/><SPLIT distance="150" swimtime="00:01:59.17"/></SPLITS></RESULT><RESULT eventid="31" heatid="340" lane="3" points="329" resultid="2533" swimtime="00:01:32.89"><SPLITS><SPLIT distance="50" swimtime="00:00:44.52"/></SPLITS></RESULT><RESULT eventid="37" heatid="406" lane="6" points="339" resultid="3028" swimtime="00:02:56.80"><SPLITS><SPLIT distance="50" swimtime="00:00:39.95"/><SPLIT distance="100" swimtime="00:01:25.57"/><SPLIT distance="150" swimtime="00:02:12.29"/></SPLITS></RESULT><RESULT eventid="39" heatid="444" lane="6" points="440" resultid="3318" swimtime="00:01:07.97"><SPLITS><SPLIT distance="50" swimtime="00:00:32.30"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="453" birthdate="2012-01-01" firstname="Greta" gender="F" lastname="Oberneder" license="458074"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="5" heatid="68" lane="1" points="359" resultid="504" swimtime="00:01:18.06"><SPLITS><SPLIT distance="50" swimtime="00:00:35.72"/></SPLITS></RESULT><RESULT eventid="11" heatid="168" lane="7" points="344" resultid="1273" swimtime="00:02:59.95"><SPLITS><SPLIT distance="50" swimtime="00:00:35.10"/><SPLIT distance="100" swimtime="00:01:22.28"/><SPLIT distance="150" swimtime="00:02:19.64"/></SPLITS></RESULT><RESULT eventid="13" heatid="202" lane="5" points="299" resultid="1532" swimtime="00:01:25.91"><SPLITS><SPLIT distance="50" swimtime="00:00:41.41"/></SPLITS></RESULT><RESULT eventid="33" heatid="359" lane="8" points="339" resultid="2674" swimtime="00:02:54.67"><SPLITS><SPLIT distance="50" swimtime="00:00:37.40"/><SPLIT distance="100" swimtime="00:01:21.25"/><SPLIT distance="150" swimtime="00:02:09.43"/></SPLITS></RESULT><RESULT eventid="35" heatid="375" lane="2" points="357" resultid="2791" swimtime="00:00:34.41"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="456" birthdate="2012-01-01" firstname="Klara" gender="F" lastname="Nagler" license="442816"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="5" heatid="68" lane="7" points="382" resultid="510" swimtime="00:01:16.46"><SPLITS><SPLIT distance="50" swimtime="00:00:35.23"/></SPLITS></RESULT><RESULT eventid="11" heatid="169" lane="1" points="404" resultid="1275" swimtime="00:02:50.55"><SPLITS><SPLIT distance="50" swimtime="00:00:36.93"/><SPLIT distance="100" swimtime="00:01:19.23"/><SPLIT distance="150" swimtime="00:02:11.68"/></SPLITS></RESULT><RESULT eventid="13" heatid="203" lane="1" points="351" resultid="1536" swimtime="00:01:21.37"><SPLITS><SPLIT distance="50" swimtime="00:00:40.29"/></SPLITS></RESULT><RESULT eventid="27" heatid="264" lane="2" points="363" resultid="1957" swimtime="00:00:37.80"><SPLITS/></RESULT><RESULT eventid="33" heatid="359" lane="6" points="376" resultid="2672" swimtime="00:02:48.75"><SPLITS><SPLIT distance="50" swimtime="00:00:36.73"/><SPLIT distance="100" swimtime="00:01:20.16"/><SPLIT distance="150" swimtime="00:02:04.60"/></SPLITS></RESULT><RESULT eventid="35" heatid="375" lane="1" points="348" resultid="2790" swimtime="00:00:34.71"><SPLITS/></RESULT><RESULT eventid="41" heatid="477" lane="7" points="395" resultid="3569" swimtime="00:06:02.77"><SPLITS><SPLIT distance="50" swimtime="00:00:38.00"/><SPLIT distance="100" swimtime="00:01:23.57"/><SPLIT distance="150" swimtime="00:02:09.42"/><SPLIT distance="200" swimtime="00:02:55.75"/><SPLIT distance="250" swimtime="00:03:47.33"/><SPLIT distance="300" swimtime="00:04:40.69"/><SPLIT distance="350" swimtime="00:05:22.73"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="464" birthdate="2006-01-01" firstname="Lena" gender="F" lastname="Gerl" license="370044"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="5" heatid="71" lane="4" points="593" resultid="531" swimtime="00:01:06.01"><SPLITS><SPLIT distance="50" swimtime="00:00:30.09"/></SPLITS></RESULT><RESULT eventid="9" heatid="131" lane="3" points="612" resultid="992" swimtime="00:00:27.87"><SPLITS/></RESULT><RESULT eventid="29" heatid="307" lane="4" points="632" resultid="2286" swimtime="00:02:11.61"><SPLITS><SPLIT distance="50" swimtime="00:00:30.10"/><SPLIT distance="100" swimtime="00:01:03.94"/><SPLIT distance="150" swimtime="00:01:38.08"/></SPLITS></RESULT><RESULT eventid="35" heatid="382" lane="3" points="542" resultid="2846" swimtime="00:00:29.96"><SPLITS/></RESULT><RESULT eventid="39" heatid="450" lane="4" points="649" resultid="3361" swimtime="00:00:59.71"><SPLITS><SPLIT distance="50" swimtime="00:00:28.57"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="468" birthdate="2014-01-01" firstname="Alexander" gender="M" lastname="Mamatov" license="449264"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="6" heatid="72" lane="1" points="146" resultid="536" swimtime="00:01:33.83"><SPLITS><SPLIT distance="50" swimtime="00:00:41.00"/></SPLITS></RESULT><RESULT eventid="8" heatid="95" lane="3" points="215" resultid="714" swimtime="00:03:30.20"><SPLITS><SPLIT distance="50" swimtime="00:00:49.10"/><SPLIT distance="100" swimtime="00:01:42.16"/><SPLIT distance="150" swimtime="00:02:38.18"/></SPLITS></RESULT><RESULT eventid="10" heatid="141" lane="8" points="196" resultid="1066" swimtime="00:00:35.95"><SPLITS/></RESULT><RESULT eventid="12" heatid="179" lane="3" points="234" resultid="1352" swimtime="00:03:04.99"><SPLITS><SPLIT distance="50" swimtime="00:00:42.07"/><SPLIT distance="100" swimtime="00:01:29.55"/><SPLIT distance="150" swimtime="00:02:25.01"/></SPLITS></RESULT><RESULT eventid="24" heatid="245" lane="5" resultid="1824" swimtime="00:00:49.20"><SPLITS/></RESULT><RESULT eventid="30" heatid="317" lane="5" points="251" resultid="2362" swimtime="00:02:41.49"><SPLITS><SPLIT distance="50" swimtime="00:00:36.11"/><SPLIT distance="100" swimtime="00:01:17.14"/><SPLIT distance="150" swimtime="00:01:59.73"/></SPLITS></RESULT><RESULT eventid="32" heatid="350" lane="8" points="195" resultid="2611" swimtime="00:01:38.07"><SPLITS><SPLIT distance="50" swimtime="00:00:46.18"/></SPLITS></RESULT><RESULT eventid="36" heatid="389" lane="8" points="145" resultid="2901" swimtime="00:00:42.35"><SPLITS/></RESULT><RESULT eventid="40" heatid="462" lane="7" points="242" resultid="3458" swimtime="00:01:15.15"><SPLITS><SPLIT distance="50" swimtime="00:00:35.32"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="469" birthdate="2014-01-01" firstname="Niklas" gender="M" lastname="Markgraf" license="449254"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="6" heatid="72" lane="2" points="170" resultid="537" swimtime="00:01:29.18"><SPLITS><SPLIT distance="50" swimtime="00:00:40.55"/></SPLITS></RESULT><RESULT eventid="10" heatid="141" lane="2" points="253" resultid="1060" swimtime="00:00:33.03"><SPLITS/></RESULT><RESULT eventid="12" heatid="180" lane="3" points="244" resultid="1360" swimtime="00:03:02.38"><SPLITS><SPLIT distance="50" swimtime="00:00:39.28"/><SPLIT distance="100" swimtime="00:01:27.17"/><SPLIT distance="150" swimtime="00:02:23.34"/></SPLITS></RESULT><RESULT eventid="14" heatid="220" lane="1" points="197" resultid="1667" swimtime="00:01:28.59"><SPLITS><SPLIT distance="50" swimtime="00:00:45.44"/></SPLITS></RESULT><RESULT eventid="20" heatid="236" lane="5" resultid="1773" swimtime="00:00:51.74"><SPLITS/></RESULT><RESULT eventid="28" heatid="280" lane="7" points="196" resultid="2083" swimtime="00:00:40.75"><SPLITS/></RESULT><RESULT eventid="30" heatid="317" lane="1" points="230" resultid="2358" swimtime="00:02:46.27"><SPLITS><SPLIT distance="50" swimtime="00:00:37.89"/><SPLIT distance="100" swimtime="00:01:21.78"/><SPLIT distance="150" swimtime="00:02:05.12"/></SPLITS></RESULT><RESULT eventid="38" heatid="416" lane="5" points="210" resultid="3103" swimtime="00:03:08.26"><SPLITS><SPLIT distance="50" swimtime="00:00:44.34"/><SPLIT distance="100" swimtime="00:01:31.62"/><SPLIT distance="150" swimtime="00:02:21.98"/></SPLITS></RESULT><RESULT eventid="40" heatid="462" lane="6" points="270" resultid="3457" swimtime="00:01:12.45"><SPLITS><SPLIT distance="50" swimtime="00:00:34.47"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="471" birthdate="2013-01-01" firstname="Anton" gender="M" lastname="Hubert" license="443842"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="6" heatid="72" lane="7" points="112" resultid="542" swimtime="00:01:42.40"><SPLITS><SPLIT distance="50" swimtime="00:00:46.34"/></SPLITS></RESULT><RESULT eventid="8" heatid="95" lane="2" points="223" resultid="713" swimtime="00:03:27.59"><SPLITS><SPLIT distance="50" swimtime="00:00:49.79"/><SPLIT distance="100" swimtime="00:01:42.21"/><SPLIT distance="150" swimtime="00:02:39.08"/></SPLITS></RESULT><RESULT eventid="10" heatid="142" lane="7" points="209" resultid="1073" swimtime="00:00:35.23"><SPLITS/></RESULT><RESULT eventid="14" heatid="219" lane="4" points="192" resultid="1662" swimtime="00:01:29.39"><SPLITS><SPLIT distance="50" swimtime="00:00:42.72"/></SPLITS></RESULT><RESULT eventid="28" heatid="281" lane="3" points="178" resultid="2087" swimtime="00:00:42.12"><SPLITS/></RESULT><RESULT eventid="30" heatid="316" lane="2" points="211" resultid="2351" swimtime="00:02:51.26"><SPLITS><SPLIT distance="50" swimtime="00:00:39.70"/><SPLIT distance="100" swimtime="00:01:24.27"/><SPLIT distance="150" swimtime="00:02:10.11"/></SPLITS></RESULT><RESULT eventid="38" heatid="416" lane="3" points="209" resultid="3101" swimtime="00:03:08.42"><SPLITS><SPLIT distance="50" swimtime="00:00:46.69"/><SPLIT distance="100" swimtime="00:01:34.55"/><SPLIT distance="150" swimtime="00:02:23.72"/></SPLITS></RESULT><RESULT eventid="40" heatid="461" lane="5" points="178" resultid="3448" swimtime="00:01:23.22"><SPLITS><SPLIT distance="50" swimtime="00:00:39.69"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="478" birthdate="2013-01-01" firstname="Alexander" gender="M" lastname="Hutchinson Riquelme" license="443849"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="6" heatid="75" lane="1" points="234" resultid="559" swimtime="00:01:20.17"><SPLITS><SPLIT distance="50" swimtime="00:00:39.09"/></SPLITS></RESULT><RESULT eventid="8" heatid="97" lane="8" points="226" resultid="733" swimtime="00:03:26.51"><SPLITS><SPLIT distance="50" swimtime="00:00:48.69"/><SPLIT distance="100" swimtime="00:01:41.89"/><SPLIT distance="150" swimtime="00:02:35.97"/></SPLITS></RESULT><RESULT eventid="10" heatid="142" lane="5" points="221" resultid="1071" swimtime="00:00:34.56"><SPLITS/></RESULT><RESULT eventid="12" heatid="181" lane="2" points="260" resultid="1367" swimtime="00:02:58.61"><SPLITS><SPLIT distance="50" swimtime="00:00:37.22"/><SPLIT distance="100" swimtime="00:01:26.44"/><SPLIT distance="150" swimtime="00:02:20.80"/></SPLITS></RESULT><RESULT eventid="22" heatid="239" lane="4" resultid="1787" swimtime="00:00:51.03"><SPLITS/></RESULT><RESULT eventid="28" heatid="280" lane="2" points="183" resultid="2078" swimtime="00:00:41.71"><SPLITS/></RESULT><RESULT eventid="30" heatid="317" lane="3" points="251" resultid="2360" swimtime="00:02:41.56"><SPLITS><SPLIT distance="50" swimtime="00:00:37.32"/><SPLIT distance="100" swimtime="00:01:19.44"/><SPLIT distance="150" swimtime="00:02:02.85"/></SPLITS></RESULT><RESULT eventid="36" heatid="391" lane="8" points="251" resultid="2917" swimtime="00:00:35.26"><SPLITS/></RESULT><RESULT eventid="40" heatid="462" lane="3" points="252" resultid="3454" swimtime="00:01:14.14"><SPLITS><SPLIT distance="50" swimtime="00:00:36.35"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="483" birthdate="2012-01-01" firstname="Luis" gender="M" lastname="Ewald" license="442810"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="6" heatid="76" lane="1" points="307" resultid="567" swimtime="00:01:13.27"><SPLITS><SPLIT distance="50" swimtime="00:00:34.76"/></SPLITS></RESULT><RESULT eventid="8" heatid="99" lane="2" points="353" resultid="742" swimtime="00:02:58.20"><SPLITS><SPLIT distance="50" swimtime="00:00:41.64"/><SPLIT distance="100" swimtime="00:01:27.00"/><SPLIT distance="150" swimtime="00:02:13.40"/></SPLITS></RESULT><RESULT eventid="12" heatid="185" lane="5" points="350" resultid="1400" swimtime="00:02:41.62"><SPLITS><SPLIT distance="50" swimtime="00:00:34.77"/><SPLIT distance="100" swimtime="00:01:18.26"/><SPLIT distance="150" swimtime="00:02:05.46"/></SPLITS></RESULT><RESULT eventid="34" heatid="361" lane="5" points="284" resultid="2686" swimtime="00:02:47.71"><SPLITS><SPLIT distance="50" swimtime="00:00:35.05"/><SPLIT distance="100" swimtime="00:01:18.32"/><SPLIT distance="150" swimtime="00:02:02.79"/></SPLITS></RESULT><RESULT eventid="36" heatid="394" lane="8" points="305" resultid="2941" swimtime="00:00:33.08"><SPLITS/></RESULT><RESULT eventid="38" heatid="418" lane="1" points="300" resultid="3114" swimtime="00:02:47.04"><SPLITS><SPLIT distance="50" swimtime="00:00:39.95"/><SPLIT distance="100" swimtime="00:01:22.26"/><SPLIT distance="150" swimtime="00:02:05.53"/></SPLITS></RESULT><RESULT eventid="42" heatid="479" lane="1" resultid="3578" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="486" birthdate="2010-01-01" firstname="Daniel" gender="M" lastname="Gross" license="415119"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="6" heatid="76" lane="6" points="310" resultid="572" swimtime="00:01:13.00"><SPLITS><SPLIT distance="50" swimtime="00:00:31.69"/></SPLITS></RESULT><RESULT eventid="10" heatid="150" lane="5" points="415" resultid="1134" swimtime="00:00:28.02"><SPLITS/></RESULT><RESULT eventid="30" heatid="322" lane="4" points="429" resultid="2399" swimtime="00:02:15.14"><SPLITS><SPLIT distance="50" swimtime="00:00:30.40"/><SPLIT distance="100" swimtime="00:01:04.52"/><SPLIT distance="150" swimtime="00:01:39.54"/></SPLITS></RESULT><RESULT eventid="36" heatid="395" lane="8" points="336" resultid="2949" swimtime="00:00:32.03"><SPLITS/></RESULT><RESULT eventid="40" heatid="470" lane="2" points="449" resultid="3515" swimtime="00:01:01.16"><SPLITS><SPLIT distance="50" swimtime="00:00:28.99"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="498" birthdate="2006-01-01" firstname="Nico" gender="M" lastname="Stuber" license="347959"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="6" heatid="79" lane="2" points="450" resultid="591" swimtime="00:01:04.50"><SPLITS><SPLIT distance="50" swimtime="00:00:28.59"/></SPLITS></RESULT><RESULT eventid="10" heatid="156" lane="8" points="453" resultid="1183" swimtime="00:00:27.21"><SPLITS/></RESULT><RESULT eventid="14" heatid="225" lane="8" points="408" resultid="1711" swimtime="00:01:09.55"><SPLITS><SPLIT distance="50" swimtime="00:00:33.67"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="501" birthdate="2008-01-01" firstname="David" gender="M" lastname="Cicero" license="412141"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="6" heatid="80" lane="4" points="536" resultid="600" swimtime="00:01:00.87"><SPLITS><SPLIT distance="50" swimtime="00:00:28.00"/></SPLITS></RESULT><RESULT eventid="10" heatid="157" lane="7" points="602" resultid="1190" swimtime="00:00:24.76"><SPLITS/></RESULT><RESULT eventid="14" heatid="225" lane="4" points="626" resultid="1707" swimtime="00:01:00.29"><SPLITS><SPLIT distance="50" swimtime="00:00:28.61"/></SPLITS></RESULT><RESULT eventid="28" heatid="287" lane="4" points="630" resultid="2135" swimtime="00:00:27.65"><SPLITS/></RESULT><RESULT eventid="36" heatid="400" lane="5" points="571" resultid="2985" swimtime="00:00:26.84"><SPLITS/></RESULT><RESULT eventid="38" heatid="419" lane="4" points="573" resultid="3122" swimtime="00:02:14.70"><SPLITS><SPLIT distance="50" swimtime="00:00:30.66"/><SPLIT distance="100" swimtime="00:01:05.30"/><SPLIT distance="150" swimtime="00:01:40.34"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="529" birthdate="2011-01-01" firstname="Maya Zoe" gender="F" lastname="Orth" license="424437"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="9" heatid="128" lane="5" points="456" resultid="971" swimtime="00:00:30.74"><SPLITS/></RESULT><RESULT eventid="13" heatid="206" lane="1" points="334" resultid="1560" swimtime="00:01:22.73"><SPLITS><SPLIT distance="50" swimtime="00:00:40.82"/></SPLITS></RESULT><RESULT eventid="27" heatid="269" lane="1" points="394" resultid="1996" swimtime="00:00:36.80"><SPLITS/></RESULT><RESULT eventid="29" heatid="304" lane="7" points="420" resultid="2267" swimtime="00:02:30.76"><SPLITS><SPLIT distance="50" swimtime="00:00:34.07"/><SPLIT distance="100" swimtime="00:01:13.40"/><SPLIT distance="150" swimtime="00:01:52.79"/></SPLITS></RESULT><RESULT eventid="37" heatid="408" lane="3" points="359" resultid="3041" swimtime="00:02:53.46"><SPLITS><SPLIT distance="50" swimtime="00:00:40.52"/><SPLIT distance="100" swimtime="00:01:24.83"/><SPLIT distance="150" swimtime="00:02:09.53"/></SPLITS></RESULT><RESULT eventid="39" heatid="447" lane="2" points="441" resultid="3337" swimtime="00:01:07.93"><SPLITS><SPLIT distance="50" swimtime="00:00:32.62"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="536" birthdate="2012-01-01" firstname="Eric-Teodor" gender="M" lastname="Mantali" license="498665"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="10" heatid="132" lane="4" resultid="998" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="30" heatid="308" lane="6" points="117" resultid="2295" swimtime="00:03:28.31"><SPLITS><SPLIT distance="50" swimtime="00:00:42.93"/><SPLIT distance="100" swimtime="00:01:35.78"/><SPLIT distance="150" swimtime="00:02:33.50"/></SPLITS></RESULT><RESULT eventid="40" heatid="451" lane="7" points="128" resultid="3372" swimtime="00:01:32.85"><SPLITS><SPLIT distance="50" swimtime="00:00:42.12"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="545" birthdate="2014-01-01" firstname="Daniel" gender="M" lastname="Löw" license="449263"><HANDICAP/><ENTRIES/><RESULTS><RESULT comment="14:43 Start vor dem Startsignal" eventid="10" heatid="140" lane="2" resultid="1053" status="DSQ" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="14" heatid="218" lane="1" points="178" resultid="1651" swimtime="00:01:31.67"><SPLITS><SPLIT distance="50" swimtime="00:00:47.13"/></SPLITS></RESULT><RESULT eventid="28" heatid="279" lane="5" points="167" resultid="2073" swimtime="00:00:43.03"><SPLITS/></RESULT><RESULT eventid="30" heatid="311" lane="4" points="161" resultid="2315" swimtime="00:03:07.42"><SPLITS><SPLIT distance="50" swimtime="00:00:42.36"/><SPLIT distance="100" swimtime="00:01:31.50"/><SPLIT distance="150" swimtime="00:02:20.98"/></SPLITS></RESULT><RESULT eventid="38" heatid="415" lane="5" points="182" resultid="3095" swimtime="00:03:17.15"><SPLITS><SPLIT distance="50" swimtime="00:00:49.82"/><SPLIT distance="100" swimtime="00:01:40.39"/><SPLIT distance="150" swimtime="00:02:31.12"/></SPLITS></RESULT><RESULT eventid="40" heatid="458" lane="7" points="155" resultid="3427" swimtime="00:01:27.11"><SPLITS><SPLIT distance="50" swimtime="00:00:42.18"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="566" birthdate="2015-01-01" firstname="Maximilian" gender="M" lastname="Rottmair" license="482345"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="14" heatid="210" lane="8" resultid="1597" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="28" heatid="273" lane="3" resultid="2026" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="30" heatid="308" lane="5" resultid="2294" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="40" heatid="451" lane="2" resultid="3367" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="567" birthdate="2014-01-01" firstname="Maximilian" gender="M" lastname="Findel" license="449253"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="14" heatid="211" lane="2" resultid="1599" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="28" heatid="276" lane="6" points="130" resultid="2052" swimtime="00:00:46.78"><SPLITS/></RESULT><RESULT eventid="30" heatid="309" lane="8" points="102" resultid="2303" swimtime="00:03:38.00"><SPLITS><SPLIT distance="50" swimtime="00:00:50.20"/><SPLIT distance="100" swimtime="00:01:48.30"/><SPLIT distance="150" swimtime="00:02:49.73"/></SPLITS></RESULT><RESULT eventid="40" heatid="453" lane="5" points="99" resultid="3386" swimtime="00:01:41.03"><SPLITS><SPLIT distance="50" swimtime="00:00:47.79"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="573" birthdate="2015-01-01" firstname="Zoe" gender="F" lastname="Vout" license="471995"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="27" heatid="255" lane="1" points="116" resultid="1884" swimtime="00:00:55.18"><SPLITS/></RESULT><RESULT eventid="31" heatid="327" lane="6" points="105" resultid="2433" swimtime="00:02:15.86"><SPLITS><SPLIT distance="50" swimtime="00:01:02.12"/></SPLITS></RESULT><RESULT eventid="37" heatid="401" lane="3" points="119" resultid="2989" swimtime="00:04:10.70"><SPLITS><SPLIT distance="50" swimtime="00:00:57.25"/><SPLIT distance="100" swimtime="00:02:02.92"/><SPLIT distance="150" swimtime="00:03:08.74"/></SPLITS></RESULT><RESULT eventid="39" heatid="420" lane="5" points="105" resultid="3129" swimtime="00:01:49.55"><SPLITS><SPLIT distance="50" swimtime="00:00:51.99"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="576" birthdate="2015-01-01" firstname="Milana" gender="F" lastname="Schneider" license="471996"><HANDICAP/><ENTRIES/><RESULTS><RESULT comment="09:10 Start vor dem Startsignal" eventid="27" heatid="257" lane="1" resultid="1900" status="DSQ" swimtime="NT"><SPLITS/></RESULT><RESULT comment="12:01 Start vor dem Startsignal" eventid="31" heatid="329" lane="3" resultid="2445" status="DSQ" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="39" heatid="424" lane="7" points="118" resultid="3161" swimtime="00:01:45.15"><SPLITS><SPLIT distance="50" swimtime="00:00:46.39"/></SPLITS></RESULT></RESULTS></ATHLETE></ATHLETES><RELAYS/></CLUB><CLUB code="4330" name="SSG Neptun Germering" nation="GER" region="02" shortname="Germerng" type="CLUB"><CONTACT city="Germering" email="gabisommer64@gmail.com" name="Sommer, Gabi" phone="089-8405373" street="Kerschensteinerstraße 94" zip="82110"/><OFFICIALS/><ATHLETES><ATHLETE athleteid="47" birthdate="2015-01-01" firstname="Alicia" gender="F" lastname="Dizerens" license="465334"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="7" lane="3" points="156" resultid="47" swimtime="00:00:54.35"><SPLITS/></RESULT><RESULT eventid="9" heatid="112" lane="4" points="211" resultid="844" swimtime="00:00:39.74"><SPLITS/></RESULT><RESULT eventid="13" heatid="195" lane="7" points="165" resultid="1478" swimtime="00:01:44.56"><SPLITS><SPLIT distance="50" swimtime="00:00:49.40"/></SPLITS></RESULT><RESULT eventid="27" heatid="260" lane="4" points="193" resultid="1927" swimtime="00:00:46.61"><SPLITS/></RESULT><RESULT eventid="29" heatid="291" lane="4" points="165" resultid="2161" swimtime="00:03:25.79"><SPLITS><SPLIT distance="50" swimtime="00:00:44.62"/><SPLIT distance="100" swimtime="00:01:38.06"/><SPLIT distance="150" swimtime="00:02:33.51"/></SPLITS></RESULT><RESULT eventid="35" heatid="364" lane="4" points="67" resultid="2706" swimtime="00:01:00.12"><SPLITS/></RESULT><RESULT eventid="39" heatid="428" lane="7" points="156" resultid="3192" swimtime="00:01:36.00"><SPLITS><SPLIT distance="50" swimtime="00:00:44.32"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="61" birthdate="2015-01-01" firstname="Malia" gender="F" lastname="Link" license="463804"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="9" lane="1" points="179" resultid="61" swimtime="00:00:51.90"><SPLITS/></RESULT><RESULT eventid="9" heatid="111" lane="5" points="187" resultid="837" swimtime="00:00:41.35"><SPLITS/></RESULT><RESULT eventid="13" heatid="195" lane="3" points="151" resultid="1474" swimtime="00:01:47.73"><SPLITS><SPLIT distance="50" swimtime="00:00:52.14"/></SPLITS></RESULT><RESULT eventid="27" heatid="260" lane="6" points="165" resultid="1929" swimtime="00:00:49.18"><SPLITS/></RESULT><RESULT eventid="31" heatid="332" lane="1" points="175" resultid="2467" swimtime="00:01:54.52"><SPLITS><SPLIT distance="50" swimtime="00:00:55.59"/></SPLITS></RESULT><RESULT eventid="39" heatid="427" lane="3" points="170" resultid="3180" swimtime="00:01:33.32"><SPLITS><SPLIT distance="50" swimtime="00:00:43.83"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="106" birthdate="2014-01-01" firstname="Nora" gender="F" lastname="Imaschewski" license="449497"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="14" lane="6" points="210" resultid="106" swimtime="00:00:49.29"><SPLITS/></RESULT><RESULT eventid="7" heatid="85" lane="8" points="211" resultid="640" swimtime="00:03:53.16"><SPLITS><SPLIT distance="50" swimtime="00:00:53.72"/><SPLIT distance="100" swimtime="00:01:52.08"/><SPLIT distance="150" swimtime="00:02:54.67"/></SPLITS></RESULT><RESULT eventid="9" heatid="111" lane="7" points="224" resultid="839" swimtime="00:00:38.93"><SPLITS/></RESULT><RESULT eventid="13" heatid="197" lane="8" points="181" resultid="1495" swimtime="00:01:41.53"><SPLITS><SPLIT distance="50" swimtime="00:00:50.03"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="113" birthdate="2011-01-01" firstname="Lara" gender="F" lastname="Dizerens" license="438350"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="15" lane="5" points="271" resultid="113" swimtime="00:00:45.25"><SPLITS/></RESULT><RESULT eventid="5" heatid="64" lane="7" points="185" resultid="479" swimtime="00:01:37.29"><SPLITS><SPLIT distance="50" swimtime="00:00:40.45"/></SPLITS></RESULT><RESULT eventid="9" heatid="117" lane="7" points="381" resultid="886" swimtime="00:00:32.65"><SPLITS/></RESULT><RESULT eventid="11" heatid="160" lane="5" points="279" resultid="1207" swimtime="00:03:12.94"><SPLITS><SPLIT distance="50" swimtime="00:00:38.96"/><SPLIT distance="100" swimtime="00:01:30.15"/><SPLIT distance="150" swimtime="00:02:25.56"/></SPLITS></RESULT><RESULT eventid="27" heatid="263" lane="2" points="302" resultid="1949" swimtime="00:00:40.19"><SPLITS/></RESULT><RESULT eventid="29" heatid="292" lane="8" points="265" resultid="2173" swimtime="00:02:55.77"><SPLITS><SPLIT distance="50" swimtime="00:00:41.71"/><SPLIT distance="100" swimtime="00:01:27.56"/><SPLIT distance="150" swimtime="00:02:15.62"/></SPLITS></RESULT><RESULT eventid="35" heatid="371" lane="3" points="279" resultid="2761" swimtime="00:00:37.37"><SPLITS/></RESULT><RESULT eventid="39" heatid="432" lane="8" points="320" resultid="3225" swimtime="00:01:15.53"><SPLITS><SPLIT distance="50" swimtime="00:00:37.37"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="145" birthdate="2011-01-01" firstname="Annika" gender="F" lastname="Arnold" license="438132"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="19" lane="5" points="393" resultid="145" swimtime="00:00:40.00"><SPLITS/></RESULT><RESULT eventid="3" heatid="46" lane="1" points="323" resultid="344" swimtime="00:05:44.53"><SPLITS><SPLIT distance="100" swimtime="00:01:31.78"/><SPLIT distance="200" swimtime="00:02:48.84"/><SPLIT distance="300" swimtime="00:04:18.59"/></SPLITS></RESULT><RESULT eventid="9" heatid="121" lane="2" points="367" resultid="913" swimtime="00:00:33.04"><SPLITS/></RESULT><RESULT eventid="27" heatid="263" lane="6" points="314" resultid="1953" swimtime="00:00:39.68"><SPLITS/></RESULT><RESULT eventid="39" heatid="441" lane="2" points="370" resultid="3290" swimtime="00:01:11.98"><SPLITS><SPLIT distance="50" swimtime="00:00:34.56"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="152" birthdate="2006-01-01" firstname="Vanessa" gender="F" lastname="Golda" license="365915"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="20" lane="4" points="403" resultid="152" swimtime="00:00:39.66"><SPLITS/></RESULT><RESULT eventid="7" heatid="89" lane="2" points="345" resultid="666" swimtime="00:03:18.04"><SPLITS><SPLIT distance="50" swimtime="00:00:44.44"/><SPLIT distance="100" swimtime="00:01:33.97"/><SPLIT distance="150" swimtime="00:02:25.37"/></SPLITS></RESULT><RESULT eventid="9" heatid="125" lane="6" points="466" resultid="949" swimtime="00:00:30.52"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="158" birthdate="2011-01-01" firstname="Antonia" gender="F" lastname="Jost" license="451122"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="21" lane="2" points="437" resultid="158" swimtime="00:00:38.61"><SPLITS/></RESULT><RESULT eventid="3" heatid="46" lane="3" points="333" resultid="346" swimtime="00:05:40.78"><SPLITS><SPLIT distance="100" swimtime="00:01:19.36"/><SPLIT distance="200" swimtime="00:02:47.81"/><SPLIT distance="300" swimtime="00:04:17.04"/></SPLITS></RESULT><RESULT eventid="9" heatid="126" lane="8" points="456" resultid="958" swimtime="00:00:30.74"><SPLITS/></RESULT><RESULT eventid="29" heatid="302" lane="4" points="396" resultid="2248" swimtime="00:02:33.84"><SPLITS><SPLIT distance="50" swimtime="00:00:35.69"/><SPLIT distance="100" swimtime="00:01:15.09"/><SPLIT distance="150" swimtime="00:01:54.86"/></SPLITS></RESULT><RESULT eventid="35" heatid="377" lane="1" points="401" resultid="2806" swimtime="00:00:33.12"><SPLITS/></RESULT><RESULT eventid="39" heatid="443" lane="2" points="444" resultid="3306" swimtime="00:01:07.76"><SPLITS><SPLIT distance="50" swimtime="00:00:33.29"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="162" birthdate="2008-01-01" firstname="Gabriela" gender="F" lastname="Rodriguez" license="488158"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="21" lane="7" resultid="162" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="9" heatid="121" lane="8" resultid="919" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="13" heatid="205" lane="2" resultid="1553" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="27" heatid="270" lane="7" resultid="2009" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="35" heatid="381" lane="8" resultid="2843" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="186" birthdate="2007-01-01" firstname="Felicitas" gender="F" lastname="Holderer" license="365916"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="24" lane="8" points="410" resultid="186" swimtime="00:00:39.42"><SPLITS/></RESULT><RESULT eventid="9" heatid="131" lane="5" points="577" resultid="993" swimtime="00:00:28.42"><SPLITS/></RESULT><RESULT eventid="11" heatid="172" lane="8" points="452" resultid="1306" swimtime="00:02:44.26"><SPLITS><SPLIT distance="50" swimtime="00:00:35.00"/><SPLIT distance="100" swimtime="00:01:20.33"/><SPLIT distance="150" swimtime="00:02:09.12"/></SPLITS></RESULT><RESULT eventid="27" heatid="270" lane="6" points="425" resultid="2008" swimtime="00:00:35.86"><SPLITS/></RESULT><RESULT eventid="31" heatid="342" lane="5" points="375" resultid="2551" swimtime="00:01:28.89"><SPLITS><SPLIT distance="50" swimtime="00:00:40.11"/></SPLITS></RESULT><RESULT eventid="35" heatid="381" lane="1" points="370" resultid="2836" swimtime="00:00:34.02"><SPLITS/></RESULT><RESULT eventid="39" heatid="450" lane="8" points="488" resultid="3365" swimtime="00:01:05.67"><SPLITS><SPLIT distance="50" swimtime="00:00:31.14"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="230" birthdate="2014-01-01" firstname="Patrick" gender="M" lastname="Calil-Hanna" license="458803"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="31" lane="2" points="130" resultid="230" swimtime="00:00:51.12"><SPLITS/></RESULT><RESULT eventid="8" heatid="94" lane="7" points="151" resultid="710" swimtime="00:03:56.24"><SPLITS><SPLIT distance="50" swimtime="00:00:52.38"/><SPLIT distance="100" swimtime="00:01:53.96"/><SPLIT distance="150" swimtime="00:02:55.95"/></SPLITS></RESULT><RESULT eventid="10" heatid="137" lane="4" points="114" resultid="1032" swimtime="00:00:43.08"><SPLITS/></RESULT><RESULT eventid="14" heatid="215" lane="5" points="113" resultid="1631" swimtime="00:01:46.48"><SPLITS><SPLIT distance="50" swimtime="00:00:52.58"/></SPLITS></RESULT><RESULT eventid="28" heatid="278" lane="7" points="118" resultid="2067" swimtime="00:00:48.25"><SPLITS/></RESULT><RESULT eventid="32" heatid="347" lane="3" points="121" resultid="2584" swimtime="00:01:54.74"><SPLITS><SPLIT distance="50" swimtime="00:00:55.94"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="231" birthdate="2016-01-01" firstname="Hector" gender="M" lastname="Seemann" license="473757"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="31" lane="3" points="122" resultid="231" swimtime="00:00:52.30"><SPLITS/></RESULT><RESULT eventid="10" heatid="139" lane="5" points="151" resultid="1048" swimtime="00:00:39.23"><SPLITS/></RESULT><RESULT eventid="14" heatid="217" lane="8" points="144" resultid="1650" swimtime="00:01:38.32"><SPLITS><SPLIT distance="50" swimtime="00:00:47.24"/></SPLITS></RESULT><RESULT eventid="30" heatid="313" lane="8" points="167" resultid="2333" swimtime="00:03:05.02"><SPLITS><SPLIT distance="50" swimtime="00:00:43.33"/><SPLIT distance="100" swimtime="00:01:31.75"/><SPLIT distance="150" swimtime="00:02:20.66"/></SPLITS></RESULT><RESULT eventid="38" heatid="414" lane="6" points="161" resultid="3088" swimtime="00:03:25.48"><SPLITS><SPLIT distance="50" swimtime="00:00:48.52"/><SPLIT distance="100" swimtime="00:01:41.57"/><SPLIT distance="150" swimtime="00:02:35.99"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="243" birthdate="2012-01-01" firstname="Jakub" gender="M" lastname="Czyzewski" license="449131"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="32" lane="7" points="239" resultid="243" swimtime="00:00:41.80"><SPLITS/></RESULT><RESULT eventid="4" heatid="55" lane="2" points="231" resultid="411" swimtime="00:05:58.60"><SPLITS><SPLIT distance="100" swimtime="00:01:19.25"/><SPLIT distance="200" swimtime="00:02:52.35"/><SPLIT distance="300" swimtime="00:04:28.42"/></SPLITS></RESULT><RESULT eventid="10" heatid="143" lane="7" points="273" resultid="1080" swimtime="00:00:32.22"><SPLITS/></RESULT><RESULT eventid="14" heatid="218" lane="7" points="215" resultid="1657" swimtime="00:01:26.02"><SPLITS><SPLIT distance="50" swimtime="00:00:39.97"/></SPLITS></RESULT><RESULT eventid="28" heatid="280" lane="3" points="233" resultid="2079" swimtime="00:00:38.51"><SPLITS/></RESULT><RESULT eventid="36" heatid="388" lane="4" points="184" resultid="2889" swimtime="00:00:39.13"><SPLITS/></RESULT><RESULT eventid="40" heatid="460" lane="4" points="258" resultid="3439" swimtime="00:01:13.52"><SPLITS><SPLIT distance="50" swimtime="00:00:33.31"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="257" birthdate="2013-01-01" firstname="Lukas" gender="M" lastname="Deng" license="449132"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="34" lane="5" points="258" resultid="257" swimtime="00:00:40.72"><SPLITS/></RESULT><RESULT eventid="6" heatid="74" lane="8" points="244" resultid="558" swimtime="00:01:19.08"><SPLITS><SPLIT distance="50" swimtime="00:00:37.11"/></SPLITS></RESULT><RESULT eventid="8" heatid="98" lane="6" points="279" resultid="738" swimtime="00:03:12.68"><SPLITS><SPLIT distance="50" swimtime="00:00:44.65"/><SPLIT distance="100" swimtime="00:01:34.92"/><SPLIT distance="150" swimtime="00:02:23.92"/></SPLITS></RESULT><RESULT eventid="12" heatid="183" lane="1" points="320" resultid="1382" swimtime="00:02:46.63"><SPLITS><SPLIT distance="50" swimtime="00:00:36.54"/><SPLIT distance="100" swimtime="00:01:18.70"/><SPLIT distance="150" swimtime="00:02:10.33"/></SPLITS></RESULT><RESULT eventid="18" heatid="232" lane="7" points="332" resultid="1753" swimtime="00:10:52.57"><SPLITS><SPLIT distance="100" swimtime="00:01:16.99"/><SPLIT distance="200" swimtime="00:02:39.54"/><SPLIT distance="300" swimtime="00:04:02.63"/><SPLIT distance="400" swimtime="00:05:26.19"/><SPLIT distance="500" swimtime="00:06:49.76"/><SPLIT distance="600" swimtime="00:08:11.65"/><SPLIT distance="700" swimtime="00:09:33.33"/></SPLITS></RESULT><RESULT eventid="26" heatid="251" lane="5" resultid="1859" swimtime="00:00:50.74"><SPLITS/></RESULT><RESULT eventid="30" heatid="316" lane="6" points="315" resultid="2355" swimtime="00:02:29.84"><SPLITS><SPLIT distance="50" swimtime="00:00:35.35"/><SPLIT distance="100" swimtime="00:01:13.55"/><SPLIT distance="150" swimtime="00:01:51.93"/></SPLITS></RESULT><RESULT eventid="34" heatid="361" lane="1" points="228" resultid="2683" swimtime="00:03:00.59"><SPLITS><SPLIT distance="50" swimtime="00:00:40.00"/><SPLIT distance="100" swimtime="00:01:27.14"/><SPLIT distance="150" swimtime="00:02:14.28"/></SPLITS></RESULT><RESULT eventid="36" heatid="389" lane="1" points="236" resultid="2894" swimtime="00:00:36.02"><SPLITS/></RESULT><RESULT eventid="42" heatid="479" lane="8" points="317" resultid="3584" swimtime="00:05:57.60"><SPLITS><SPLIT distance="50" swimtime="00:00:39.73"/><SPLIT distance="100" swimtime="00:01:27.58"/><SPLIT distance="150" swimtime="00:02:14.50"/><SPLIT distance="200" swimtime="00:02:59.46"/><SPLIT distance="250" swimtime="00:03:50.35"/><SPLIT distance="300" swimtime="00:04:39.90"/><SPLIT distance="350" swimtime="00:05:19.78"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="264" birthdate="2011-01-01" firstname="Lars" gender="M" lastname="Holderer" license="423863"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="35" lane="6" points="282" resultid="264" swimtime="00:00:39.57"><SPLITS/></RESULT><RESULT eventid="8" heatid="98" lane="7" points="271" resultid="739" swimtime="00:03:14.46"><SPLITS><SPLIT distance="50" swimtime="00:00:44.62"/><SPLIT distance="100" swimtime="00:01:35.68"/><SPLIT distance="150" swimtime="00:02:24.91"/></SPLITS></RESULT><RESULT eventid="10" heatid="146" lane="6" points="298" resultid="1103" swimtime="00:00:31.29"><SPLITS/></RESULT><RESULT eventid="12" heatid="181" lane="4" points="269" resultid="1369" swimtime="00:02:56.39"><SPLITS><SPLIT distance="50" swimtime="00:00:41.10"/><SPLIT distance="100" swimtime="00:01:28.92"/><SPLIT distance="150" swimtime="00:02:16.44"/></SPLITS></RESULT><RESULT eventid="16" heatid="228" lane="6" points="295" resultid="1723" swimtime="00:21:47.87"><SPLITS><SPLIT distance="100" swimtime="00:01:17.34"/><SPLIT distance="200" swimtime="00:02:42.90"/><SPLIT distance="300" swimtime="00:04:09.69"/><SPLIT distance="400" swimtime="00:05:37.65"/><SPLIT distance="500" swimtime="00:07:05.79"/><SPLIT distance="600" swimtime="00:08:34.53"/><SPLIT distance="700" swimtime="00:10:03.03"/><SPLIT distance="800" swimtime="00:11:31.77"/><SPLIT distance="900" swimtime="00:13:00.37"/><SPLIT distance="1000" swimtime="00:14:28.23"/><SPLIT distance="1100" swimtime="00:15:56.76"/><SPLIT distance="1200" swimtime="00:17:25.07"/><SPLIT distance="1300" swimtime="00:18:54.78"/><SPLIT distance="1400" swimtime="00:20:22.38"/></SPLITS></RESULT><RESULT eventid="28" heatid="282" lane="2" points="197" resultid="2094" swimtime="00:00:40.73"><SPLITS/></RESULT><RESULT eventid="32" heatid="352" lane="8" points="247" resultid="2626" swimtime="00:01:30.61"><SPLITS><SPLIT distance="50" swimtime="00:00:43.51"/></SPLITS></RESULT><RESULT eventid="36" heatid="389" lane="5" points="161" resultid="2898" swimtime="00:00:40.87"><SPLITS/></RESULT><RESULT eventid="40" heatid="466" lane="7" points="308" resultid="3489" swimtime="00:01:09.37"><SPLITS><SPLIT distance="50" swimtime="00:00:33.22"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="273" birthdate="2011-01-01" firstname="Benjamin" gender="M" lastname="Weber" license="434655"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="36" lane="7" points="279" resultid="273" swimtime="00:00:39.68"><SPLITS/></RESULT><RESULT eventid="8" heatid="96" lane="4" points="248" resultid="721" swimtime="00:03:20.40"><SPLITS><SPLIT distance="50" swimtime="00:00:45.20"/><SPLIT distance="100" swimtime="00:01:36.87"/><SPLIT distance="150" swimtime="00:02:29.16"/></SPLITS></RESULT><RESULT eventid="10" heatid="145" lane="5" points="266" resultid="1094" swimtime="00:00:32.51"><SPLITS/></RESULT><RESULT eventid="14" heatid="220" lane="7" points="243" resultid="1672" swimtime="00:01:22.65"><SPLITS><SPLIT distance="50" swimtime="00:00:37.94"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="307" birthdate="2014-01-01" firstname="Amelie" gender="F" lastname="Schrader" license="465328"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="41" lane="2" points="168" resultid="307" swimtime="00:07:08.28"><SPLITS><SPLIT distance="100" swimtime="00:01:37.28"/><SPLIT distance="200" swimtime="00:03:26.78"/><SPLIT distance="300" swimtime="00:05:17.41"/></SPLITS></RESULT><RESULT eventid="7" heatid="85" lane="2" points="223" resultid="634" swimtime="00:03:48.87"><SPLITS><SPLIT distance="50" swimtime="00:00:51.77"/><SPLIT distance="100" swimtime="00:01:47.90"/><SPLIT distance="150" swimtime="00:02:49.74"/></SPLITS></RESULT><RESULT eventid="11" heatid="160" lane="1" points="201" resultid="1203" swimtime="00:03:35.06"><SPLITS><SPLIT distance="50" swimtime="00:00:45.27"/><SPLIT distance="100" swimtime="00:01:43.03"/><SPLIT distance="150" swimtime="00:02:46.52"/></SPLITS></RESULT><RESULT eventid="23" heatid="241" lane="3" resultid="1794" swimtime="00:00:54.33"><SPLITS/></RESULT><RESULT eventid="29" heatid="291" lane="5" points="181" resultid="2162" swimtime="00:03:19.55"><SPLITS><SPLIT distance="50" swimtime="00:00:43.30"/><SPLIT distance="100" swimtime="00:01:34.41"/><SPLIT distance="150" swimtime="00:02:29.33"/></SPLITS></RESULT><RESULT eventid="37" heatid="403" lane="5" points="178" resultid="3003" swimtime="00:03:39.21"><SPLITS><SPLIT distance="50" swimtime="00:00:51.06"/><SPLIT distance="100" swimtime="00:01:46.33"/><SPLIT distance="150" swimtime="00:02:43.88"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="308" birthdate="2013-01-01" firstname="Lou" gender="F" lastname="Wunderlich" license="465091"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="41" lane="3" points="195" resultid="308" swimtime="00:06:47.03"><SPLITS><SPLIT distance="100" swimtime="00:01:38.39"/><SPLIT distance="200" swimtime="00:03:24.50"/><SPLIT distance="300" swimtime="00:05:08.53"/></SPLITS></RESULT><RESULT comment="11:48 Start vor dem Startsignal" eventid="7" heatid="82" lane="4" resultid="613" status="DSQ" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="11" heatid="159" lane="3" points="195" resultid="1198" swimtime="00:03:37.45"><SPLITS><SPLIT distance="50" swimtime="00:00:53.15"/><SPLIT distance="100" swimtime="00:01:48.64"/><SPLIT distance="150" swimtime="00:02:50.82"/></SPLITS></RESULT><RESULT eventid="23" heatid="242" lane="2" resultid="1800" swimtime="00:00:51.56"><SPLITS/></RESULT><RESULT eventid="29" heatid="290" lane="3" points="215" resultid="2153" swimtime="00:03:08.54"><SPLITS><SPLIT distance="50" swimtime="00:00:44.85"/><SPLIT distance="100" swimtime="00:01:34.50"/><SPLIT distance="150" swimtime="00:02:23.48"/></SPLITS></RESULT><RESULT eventid="37" heatid="404" lane="3" points="181" resultid="3009" swimtime="00:03:38.03"><SPLITS><SPLIT distance="50" swimtime="00:00:53.14"/><SPLIT distance="100" swimtime="00:01:49.49"/><SPLIT distance="150" swimtime="00:02:44.71"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="309" birthdate="2013-01-01" firstname="Sophia" gender="F" lastname="Tait" license="480267"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="41" lane="4" points="190" resultid="309" swimtime="00:06:50.87"><SPLITS><SPLIT distance="100" swimtime="00:01:34.47"/><SPLIT distance="200" swimtime="00:03:21.02"/><SPLIT distance="300" swimtime="00:05:08.44"/></SPLITS></RESULT><RESULT eventid="7" heatid="86" lane="3" points="272" resultid="643" swimtime="00:03:34.38"><SPLITS><SPLIT distance="50" swimtime="00:00:48.32"/><SPLIT distance="100" swimtime="00:01:41.83"/><SPLIT distance="150" swimtime="00:02:38.70"/></SPLITS></RESULT><RESULT eventid="11" heatid="161" lane="1" points="230" resultid="1211" swimtime="00:03:25.64"><SPLITS><SPLIT distance="50" swimtime="00:00:43.44"/><SPLIT distance="100" swimtime="00:01:36.47"/><SPLIT distance="150" swimtime="00:02:35.03"/></SPLITS></RESULT><RESULT eventid="23" heatid="242" lane="8" resultid="1806" swimtime="00:00:59.82"><SPLITS/></RESULT><RESULT eventid="29" heatid="292" lane="3" points="193" resultid="2168" swimtime="00:03:15.24"><SPLITS><SPLIT distance="50" swimtime="00:00:42.98"/><SPLIT distance="100" swimtime="00:01:32.63"/><SPLIT distance="150" swimtime="00:02:26.19"/></SPLITS></RESULT><RESULT eventid="37" heatid="404" lane="7" points="204" resultid="3013" swimtime="00:03:29.23"><SPLITS><SPLIT distance="50" swimtime="00:00:46.30"/><SPLIT distance="100" swimtime="00:01:41.12"/><SPLIT distance="150" swimtime="00:02:36.00"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="310" birthdate="2013-01-01" firstname="Luisa" gender="F" lastname="Feuerhak" license="444792"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="41" lane="6" points="170" resultid="310" swimtime="00:07:06.69"><SPLITS><SPLIT distance="100" swimtime="00:01:35.66"/><SPLIT distance="200" swimtime="00:03:23.94"/><SPLIT distance="300" swimtime="00:05:16.22"/></SPLITS></RESULT><RESULT eventid="7" heatid="86" lane="6" points="262" resultid="646" swimtime="00:03:37.07"><SPLITS><SPLIT distance="50" swimtime="00:00:52.40"/><SPLIT distance="100" swimtime="00:01:49.38"/><SPLIT distance="150" swimtime="00:02:42.79"/></SPLITS></RESULT><RESULT eventid="11" heatid="159" lane="5" points="195" resultid="1200" swimtime="00:03:37.31"><SPLITS><SPLIT distance="50" swimtime="00:00:46.85"/><SPLIT distance="100" swimtime="00:01:46.73"/><SPLIT distance="150" swimtime="00:02:46.91"/></SPLITS></RESULT><RESULT eventid="23" heatid="241" lane="5" resultid="1796" swimtime="00:00:58.31"><SPLITS/></RESULT><RESULT eventid="29" heatid="291" lane="2" points="192" resultid="2159" swimtime="00:03:15.71"><SPLITS><SPLIT distance="50" swimtime="00:00:44.30"/><SPLIT distance="100" swimtime="00:01:33.98"/><SPLIT distance="150" swimtime="00:02:25.71"/></SPLITS></RESULT><RESULT eventid="37" heatid="404" lane="5" points="207" resultid="3011" swimtime="00:03:28.23"><SPLITS><SPLIT distance="50" swimtime="00:00:53.59"/><SPLIT distance="100" swimtime="00:01:47.05"/><SPLIT distance="150" swimtime="00:02:40.05"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="326" birthdate="2013-01-01" firstname="Luana Nina" gender="F" lastname="Link" license="444793"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="44" lane="5" points="243" resultid="332" swimtime="00:06:18.52"><SPLITS><SPLIT distance="100" swimtime="00:01:24.50"/><SPLIT distance="200" swimtime="00:03:01.37"/><SPLIT distance="300" swimtime="00:04:40.80"/></SPLITS></RESULT><RESULT eventid="7" heatid="86" lane="1" points="199" resultid="641" swimtime="00:03:57.69"><SPLITS><SPLIT distance="50" swimtime="00:00:54.10"/><SPLIT distance="100" swimtime="00:01:55.19"/><SPLIT distance="150" swimtime="00:02:58.71"/></SPLITS></RESULT><RESULT eventid="11" heatid="161" lane="8" points="243" resultid="1218" swimtime="00:03:21.96"><SPLITS><SPLIT distance="50" swimtime="00:00:44.04"/><SPLIT distance="100" swimtime="00:01:33.98"/><SPLIT distance="150" swimtime="00:02:34.75"/></SPLITS></RESULT><RESULT eventid="23" heatid="241" lane="4" resultid="1795" swimtime="00:00:57.28"><SPLITS/></RESULT><RESULT eventid="29" heatid="295" lane="7" points="239" resultid="2196" swimtime="00:03:01.84"><SPLITS><SPLIT distance="50" swimtime="00:00:39.07"/><SPLIT distance="100" swimtime="00:01:25.94"/><SPLIT distance="150" swimtime="00:02:13.69"/></SPLITS></RESULT><RESULT eventid="37" heatid="405" lane="7" points="244" resultid="3021" swimtime="00:03:17.35"><SPLITS><SPLIT distance="50" swimtime="00:00:46.78"/><SPLIT distance="100" swimtime="00:01:37.52"/><SPLIT distance="150" swimtime="00:02:28.28"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="357" birthdate="2009-01-01" firstname="Annika" gender="F" lastname="Tischner" license="416838"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="50" lane="1" points="312" resultid="375" swimtime="00:05:48.19"><SPLITS><SPLIT distance="100" swimtime="00:01:18.98"/><SPLIT distance="200" swimtime="00:02:46.59"/><SPLIT distance="300" swimtime="00:04:17.59"/></SPLITS></RESULT><RESULT eventid="9" heatid="126" lane="6" points="461" resultid="957" swimtime="00:00:30.64"><SPLITS/></RESULT><RESULT eventid="13" heatid="205" lane="4" points="404" resultid="1555" swimtime="00:01:17.68"><SPLITS><SPLIT distance="50" swimtime="00:00:38.39"/></SPLITS></RESULT><RESULT eventid="17" heatid="231" lane="2" points="405" resultid="1741" swimtime="00:10:55.13"><SPLITS><SPLIT distance="100" swimtime="00:01:15.17"/><SPLIT distance="200" swimtime="00:02:37.65"/><SPLIT distance="300" swimtime="00:04:00.43"/><SPLIT distance="400" swimtime="00:05:23.62"/><SPLIT distance="500" swimtime="00:06:47.40"/><SPLIT distance="600" swimtime="00:08:12.38"/><SPLIT distance="700" swimtime="00:09:36.52"/></SPLITS></RESULT><RESULT eventid="27" heatid="269" lane="3" points="411" resultid="1998" swimtime="00:00:36.28"><SPLITS/></RESULT><RESULT eventid="29" heatid="304" lane="8" points="429" resultid="2268" swimtime="00:02:29.78"><SPLITS><SPLIT distance="50" swimtime="00:00:34.97"/><SPLIT distance="100" swimtime="00:01:12.65"/><SPLIT distance="150" swimtime="00:01:53.03"/></SPLITS></RESULT><RESULT eventid="37" heatid="409" lane="5" points="364" resultid="3051" swimtime="00:02:52.62"><SPLITS><SPLIT distance="50" swimtime="00:00:41.81"/><SPLIT distance="100" swimtime="00:01:26.54"/><SPLIT distance="150" swimtime="00:02:11.39"/></SPLITS></RESULT><RESULT eventid="39" heatid="446" lane="6" points="450" resultid="3333" swimtime="00:01:07.45"><SPLITS><SPLIT distance="50" swimtime="00:00:32.57"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="376" birthdate="2010-01-01" firstname="Carys" gender="F" lastname="Wagner" license="433934"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="52" lane="6" points="590" resultid="395" swimtime="00:04:41.81"><SPLITS><SPLIT distance="100" swimtime="00:01:07.34"/><SPLIT distance="200" swimtime="00:02:18.90"/><SPLIT distance="300" swimtime="00:03:30.79"/></SPLITS></RESULT><RESULT eventid="11" heatid="174" lane="6" points="592" resultid="1320" swimtime="00:02:30.12"><SPLITS><SPLIT distance="50" swimtime="00:00:32.92"/><SPLIT distance="100" swimtime="00:01:12.12"/><SPLIT distance="150" swimtime="00:01:56.32"/></SPLITS></RESULT><RESULT eventid="13" heatid="208" lane="4" points="528" resultid="1578" swimtime="00:01:11.07"><SPLITS><SPLIT distance="50" swimtime="00:00:34.14"/></SPLITS></RESULT><RESULT eventid="37" heatid="412" lane="7" points="515" resultid="3077" swimtime="00:02:33.80"><SPLITS><SPLIT distance="100" swimtime="00:01:14.14"/></SPLITS></RESULT><RESULT eventid="41" heatid="478" lane="6" points="585" resultid="3575" swimtime="00:05:18.48"><SPLITS><SPLIT distance="50" swimtime="00:00:34.03"/><SPLIT distance="100" swimtime="00:01:15.58"/><SPLIT distance="150" swimtime="00:01:57.84"/><SPLIT distance="200" swimtime="00:02:38.20"/><SPLIT distance="250" swimtime="00:03:22.77"/><SPLIT distance="300" swimtime="00:04:08.14"/><SPLIT distance="350" swimtime="00:04:43.60"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="380" birthdate="2014-01-01" firstname="Oskar" gender="M" lastname="Stubbe" license="475469"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="53" lane="4" points="164" resultid="400" swimtime="00:06:41.59"><SPLITS><SPLIT distance="200" swimtime="00:03:19.42"/><SPLIT distance="300" swimtime="00:05:03.37"/></SPLITS></RESULT><RESULT eventid="10" heatid="140" lane="5" points="171" resultid="1056" swimtime="00:00:37.64"><SPLITS/></RESULT><RESULT eventid="14" heatid="216" lane="5" points="130" resultid="1639" swimtime="00:01:41.69"><SPLITS><SPLIT distance="50" swimtime="00:00:49.86"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="384" birthdate="2015-01-01" firstname="Timo" gender="M" lastname="Deng" license="463803"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="54" lane="5" points="149" resultid="406" swimtime="00:06:54.35"><SPLITS><SPLIT distance="100" swimtime="00:01:34.31"/><SPLIT distance="200" swimtime="00:03:24.55"/><SPLIT distance="300" swimtime="00:05:09.83"/></SPLITS></RESULT><RESULT eventid="8" heatid="94" lane="5" points="153" resultid="708" swimtime="00:03:55.18"><SPLITS><SPLIT distance="50" swimtime="00:00:53.60"/><SPLIT distance="100" swimtime="00:01:57.69"/><SPLIT distance="150" swimtime="00:02:57.52"/></SPLITS></RESULT><RESULT eventid="12" heatid="177" lane="6" points="177" resultid="1340" swimtime="00:03:22.81"><SPLITS><SPLIT distance="50" swimtime="00:00:43.25"/><SPLIT distance="100" swimtime="00:01:33.67"/><SPLIT distance="150" swimtime="00:02:37.34"/></SPLITS></RESULT><RESULT eventid="30" heatid="313" lane="2" points="154" resultid="2328" swimtime="00:03:10.07"><SPLITS><SPLIT distance="50" swimtime="00:00:41.22"/><SPLIT distance="100" swimtime="00:01:31.17"/><SPLIT distance="150" swimtime="00:02:25.47"/></SPLITS></RESULT><RESULT eventid="38" heatid="415" lane="8" points="165" resultid="3098" swimtime="00:03:23.88"><SPLITS><SPLIT distance="50" swimtime="00:00:48.03"/><SPLIT distance="100" swimtime="00:01:41.06"/><SPLIT distance="150" swimtime="00:02:36.23"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="387" birthdate="2015-01-01" firstname="Valentin" gender="M" lastname="Lekies" license="458874"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="54" lane="8" points="158" resultid="409" swimtime="00:06:46.28"><SPLITS><SPLIT distance="100" swimtime="00:01:34.23"/><SPLIT distance="200" swimtime="00:03:22.38"/><SPLIT distance="300" swimtime="00:05:08.41"/></SPLITS></RESULT><RESULT eventid="8" heatid="96" lane="6" points="166" resultid="723" swimtime="00:03:49.16"><SPLITS><SPLIT distance="50" swimtime="00:00:53.08"/><SPLIT distance="100" swimtime="00:01:52.65"/><SPLIT distance="150" swimtime="00:02:52.73"/></SPLITS></RESULT><RESULT eventid="12" heatid="176" lane="6" points="149" resultid="1333" swimtime="00:03:35.03"><SPLITS><SPLIT distance="50" swimtime="00:00:54.56"/><SPLIT distance="100" swimtime="00:01:52.04"/><SPLIT distance="150" swimtime="00:02:48.96"/></SPLITS></RESULT><RESULT eventid="30" heatid="313" lane="3" points="152" resultid="2329" swimtime="00:03:11.11"><SPLITS><SPLIT distance="50" swimtime="00:00:42.87"/><SPLIT distance="100" swimtime="00:01:33.45"/><SPLIT distance="150" swimtime="00:02:27.02"/></SPLITS></RESULT><RESULT eventid="38" heatid="415" lane="1" points="172" resultid="3091" swimtime="00:03:21.10"><SPLITS><SPLIT distance="100" swimtime="00:01:41.03"/><SPLIT distance="150" swimtime="00:02:34.68"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="404" birthdate="2011-01-01" firstname="Rüzgar" gender="M" lastname="Ugur" license="461737"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="57" lane="5" points="265" resultid="430" swimtime="00:05:42.41"><SPLITS><SPLIT distance="100" swimtime="00:01:12.59"/><SPLIT distance="200" swimtime="00:02:42.02"/><SPLIT distance="300" swimtime="00:04:13.98"/></SPLITS></RESULT><RESULT eventid="10" heatid="148" lane="5" points="383" resultid="1118" swimtime="00:00:28.78"><SPLITS/></RESULT><RESULT eventid="12" heatid="182" lane="2" points="296" resultid="1375" swimtime="00:02:51.02"><SPLITS><SPLIT distance="50" swimtime="00:00:36.10"/><SPLIT distance="100" swimtime="00:01:20.04"/><SPLIT distance="150" swimtime="00:02:13.51"/></SPLITS></RESULT><RESULT eventid="32" heatid="351" lane="5" points="269" resultid="2616" swimtime="00:01:28.04"><SPLITS><SPLIT distance="50" swimtime="00:00:39.96"/></SPLITS></RESULT><RESULT eventid="36" heatid="393" lane="7" points="317" resultid="2932" swimtime="00:00:32.66"><SPLITS/></RESULT><RESULT eventid="38" heatid="417" lane="2" points="293" resultid="3108" swimtime="00:02:48.34"><SPLITS><SPLIT distance="50" swimtime="00:00:37.39"/><SPLIT distance="100" swimtime="00:01:20.99"/><SPLIT distance="150" swimtime="00:02:07.31"/></SPLITS></RESULT><RESULT eventid="40" heatid="468" lane="7" points="378" resultid="3504" swimtime="00:01:04.77"><SPLITS><SPLIT distance="50" swimtime="00:00:30.08"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="488" birthdate="2009-01-01" firstname="Maximo" gender="M" lastname="Flath" license="464194"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="6" heatid="77" lane="2" points="367" resultid="576" swimtime="00:01:09.04"><SPLITS><SPLIT distance="50" swimtime="00:00:31.31"/></SPLITS></RESULT><RESULT eventid="10" heatid="149" lane="5" points="449" resultid="1126" swimtime="00:00:27.30"><SPLITS/></RESULT><RESULT eventid="14" heatid="223" lane="8" points="338" resultid="1696" swimtime="00:01:14.05"><SPLITS><SPLIT distance="50" swimtime="00:00:37.34"/></SPLITS></RESULT><RESULT eventid="28" heatid="284" lane="5" points="387" resultid="2112" swimtime="00:00:32.53"><SPLITS/></RESULT><RESULT eventid="36" heatid="395" lane="7" points="456" resultid="2948" swimtime="00:00:28.92"><SPLITS/></RESULT><RESULT eventid="40" heatid="468" lane="3" points="446" resultid="3500" swimtime="00:01:01.30"><SPLITS><SPLIT distance="50" swimtime="00:00:29.91"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="514" birthdate="2015-01-01" firstname="Romy" gender="F" lastname="Scheller" license="485979"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="9" heatid="109" lane="6" points="169" resultid="822" swimtime="00:00:42.76"><SPLITS/></RESULT><RESULT eventid="13" heatid="194" lane="4" points="136" resultid="1467" swimtime="00:01:51.67"><SPLITS><SPLIT distance="50" swimtime="00:00:55.30"/></SPLITS></RESULT><RESULT eventid="27" heatid="258" lane="2" points="160" resultid="1909" swimtime="00:00:49.64"><SPLITS/></RESULT><RESULT eventid="31" heatid="330" lane="2" points="134" resultid="2452" swimtime="00:02:05.29"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="528" birthdate="2004-01-01" firstname="Alessia" gender="F" lastname="Tammaro" license="333921"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="9" heatid="127" lane="2" points="465" resultid="960" swimtime="00:00:30.55"><SPLITS/></RESULT><RESULT eventid="13" heatid="209" lane="8" points="524" resultid="1589" swimtime="00:01:11.23"><SPLITS><SPLIT distance="50" swimtime="00:00:34.74"/></SPLITS></RESULT><RESULT eventid="27" heatid="272" lane="2" points="536" resultid="2019" swimtime="00:00:33.21"><SPLITS/></RESULT><RESULT eventid="35" heatid="380" lane="5" points="425" resultid="2832" swimtime="00:00:32.47"><SPLITS/></RESULT><RESULT eventid="39" heatid="447" lane="4" points="471" resultid="3339" swimtime="00:01:06.44"><SPLITS><SPLIT distance="50" swimtime="00:00:31.94"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="531" birthdate="2003-01-01" firstname="Claudia" gender="F" lastname="Dobmeier" license="299888"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="9" heatid="129" lane="5" points="477" resultid="979" swimtime="00:00:30.28"><SPLITS/></RESULT><RESULT eventid="13" heatid="208" lane="1" points="416" resultid="1575" swimtime="00:01:16.93"><SPLITS><SPLIT distance="50" swimtime="00:00:36.66"/></SPLITS></RESULT><RESULT eventid="27" heatid="271" lane="3" resultid="2012" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="35" heatid="378" lane="3" resultid="2814" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="39" heatid="448" lane="1" resultid="3343" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="547" birthdate="2011-01-01" firstname="Ole" gender="M" lastname="Plass" license="434296"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="10" heatid="143" lane="4" points="250" resultid="1077" swimtime="00:00:33.16"><SPLITS/></RESULT><RESULT eventid="12" heatid="178" lane="1" points="191" resultid="1343" swimtime="00:03:17.65"><SPLITS><SPLIT distance="50" swimtime="00:00:42.33"/><SPLIT distance="100" swimtime="00:01:29.79"/><SPLIT distance="150" swimtime="00:02:30.31"/></SPLITS></RESULT><RESULT eventid="14" heatid="218" lane="2" points="182" resultid="1652" swimtime="00:01:30.90"><SPLITS><SPLIT distance="50" swimtime="00:00:44.13"/></SPLITS></RESULT><RESULT eventid="30" heatid="315" lane="7" points="192" resultid="2348" swimtime="00:02:56.75"><SPLITS><SPLIT distance="50" swimtime="00:00:38.62"/><SPLIT distance="100" swimtime="00:01:23.54"/><SPLIT distance="150" swimtime="00:02:11.41"/></SPLITS></RESULT><RESULT eventid="36" heatid="388" lane="6" points="203" resultid="2891" swimtime="00:00:37.89"><SPLITS/></RESULT><RESULT eventid="40" heatid="461" lane="6" points="226" resultid="3449" swimtime="00:01:16.87"><SPLITS><SPLIT distance="50" swimtime="00:00:36.45"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="570" birthdate="2014-01-01" firstname="Felicia" gender="F" lastname="Schrader" license="465330"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="23" heatid="241" lane="6" resultid="1797" swimtime="00:00:57.76"><SPLITS/></RESULT><RESULT eventid="29" heatid="292" lane="6" points="213" resultid="2171" swimtime="00:03:09.13"><SPLITS><SPLIT distance="50" swimtime="00:00:42.63"/><SPLIT distance="100" swimtime="00:01:31.87"/><SPLIT distance="150" swimtime="00:02:23.12"/></SPLITS></RESULT><RESULT eventid="37" heatid="403" lane="2" resultid="3000" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="577" birthdate="2016-01-01" firstname="Leonie" gender="F" lastname="Henne" license="482273"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="27" heatid="257" lane="7" points="145" resultid="1906" swimtime="00:00:51.25"><SPLITS/></RESULT><RESULT eventid="31" heatid="330" lane="4" points="153" resultid="2454" swimtime="00:01:59.69"><SPLITS/></RESULT><RESULT eventid="39" heatid="425" lane="3" points="128" resultid="3165" swimtime="00:01:42.44"><SPLITS><SPLIT distance="50" swimtime="00:00:48.72"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="584" birthdate="2014-01-01" firstname="Lena" gender="F" lastname="Henne" license="463028"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="27" heatid="264" lane="8" points="254" resultid="1963" swimtime="00:00:42.58"><SPLITS/></RESULT><RESULT eventid="29" heatid="292" lane="2" points="163" resultid="2167" swimtime="00:03:26.60"><SPLITS><SPLIT distance="50" swimtime="00:00:43.13"/><SPLIT distance="100" swimtime="00:01:34.28"/><SPLIT distance="150" swimtime="00:02:30.74"/></SPLITS></RESULT><RESULT eventid="35" heatid="369" lane="7" points="185" resultid="2749" swimtime="00:00:42.81"><SPLITS/></RESULT><RESULT eventid="39" heatid="430" lane="3" points="209" resultid="3204" swimtime="00:01:27.04"><SPLITS><SPLIT distance="50" swimtime="00:00:40.46"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="594" birthdate="2012-01-01" firstname="Eddie" gender="M" lastname="Li" license="449133"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="28" heatid="279" lane="3" points="160" resultid="2071" swimtime="00:00:43.64"><SPLITS/></RESULT><RESULT eventid="30" heatid="315" lane="8" points="189" resultid="2349" swimtime="00:02:57.46"><SPLITS><SPLIT distance="50" swimtime="00:00:38.68"/><SPLIT distance="100" swimtime="00:01:24.23"/><SPLIT distance="150" swimtime="00:02:13.54"/></SPLITS></RESULT><RESULT eventid="36" heatid="387" lane="1" points="133" resultid="2879" swimtime="00:00:43.60"><SPLITS/></RESULT><RESULT eventid="40" heatid="461" lane="8" points="210" resultid="3451" swimtime="00:01:18.76"><SPLITS><SPLIT distance="50" swimtime="00:00:36.12"/></SPLITS></RESULT></RESULTS></ATHLETE></ATHLETES><RELAYS/></CLUB><CLUB code="4341" name="SV Hof" nation="GER" region="02" shortname="Hof" type="CLUB"><CONTACT city="Hof" country="GER" email="maler.reiss@t-online.de" fax="928191461" name="Reiss, Barbara" phone="09281/91109" street="Ziegeleiweg 6" zip="95032"/><OFFICIALS/><ATHLETES><ATHLETE athleteid="51" birthdate="2016-01-01" firstname="Coralie" gender="F" lastname="Münch" license="482662"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="7" lane="7" points="135" resultid="51" swimtime="00:00:57.06"><SPLITS/></RESULT><RESULT eventid="9" heatid="105" lane="4" points="148" resultid="788" swimtime="00:00:44.74"><SPLITS/></RESULT><RESULT eventid="13" heatid="192" lane="1" points="161" resultid="1448" swimtime="00:01:45.53"><SPLITS><SPLIT distance="50" swimtime="00:00:51.46"/></SPLITS></RESULT><RESULT eventid="27" heatid="257" lane="3" points="180" resultid="1902" swimtime="00:00:47.72"><SPLITS/></RESULT><RESULT eventid="31" heatid="328" lane="2" points="144" resultid="2436" swimtime="00:02:02.21"><SPLITS><SPLIT distance="50" swimtime="00:00:58.33"/></SPLITS></RESULT><RESULT comment="14:49 Die Sportlerin hat während der Schwimmstrecke ihre Bahn verlassen" eventid="37" heatid="401" lane="4" resultid="2990" status="DSQ" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="39" heatid="422" lane="7" points="114" resultid="3145" swimtime="00:01:46.55"><SPLITS><SPLIT distance="50" swimtime="00:00:49.98"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="118" birthdate="2012-01-01" firstname="Melina" gender="F" lastname="Schmidt" license="452716"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="16" lane="2" points="269" resultid="118" swimtime="00:00:45.34"><SPLITS/></RESULT><RESULT eventid="7" heatid="84" lane="7" points="259" resultid="631" swimtime="00:03:37.79"><SPLITS><SPLIT distance="50" swimtime="00:00:48.92"/><SPLIT distance="100" swimtime="00:01:45.02"/><SPLIT distance="150" swimtime="00:02:42.46"/></SPLITS></RESULT><RESULT eventid="9" heatid="113" lane="1" points="228" resultid="849" swimtime="00:00:38.69"><SPLITS/></RESULT><RESULT eventid="13" heatid="196" lane="3" points="160" resultid="1482" swimtime="00:01:45.78"><SPLITS/></RESULT><RESULT eventid="27" heatid="261" lane="8" points="198" resultid="1939" swimtime="00:00:46.22"><SPLITS/></RESULT><RESULT eventid="31" heatid="336" lane="2" points="241" resultid="2500" swimtime="00:01:43.00"><SPLITS><SPLIT distance="50" swimtime="00:00:49.09"/></SPLITS></RESULT><RESULT eventid="39" heatid="429" lane="4" points="179" resultid="3197" swimtime="00:01:31.65"><SPLITS><SPLIT distance="50" swimtime="00:00:42.33"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="131" birthdate="2010-01-01" firstname="Elodie" gender="F" lastname="Münch" license="402456"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="17" lane="7" points="267" resultid="131" swimtime="00:00:45.47"><SPLITS/></RESULT><RESULT eventid="5" heatid="65" lane="3" points="212" resultid="483" swimtime="00:01:32.96"><SPLITS><SPLIT distance="50" swimtime="00:00:41.85"/></SPLITS></RESULT><RESULT eventid="9" heatid="122" lane="1" points="377" resultid="920" swimtime="00:00:32.76"><SPLITS/></RESULT><RESULT eventid="13" heatid="203" lane="5" points="318" resultid="1540" swimtime="00:01:24.09"><SPLITS><SPLIT distance="50" swimtime="00:00:40.84"/></SPLITS></RESULT><RESULT eventid="27" heatid="266" lane="6" points="322" resultid="1977" swimtime="00:00:39.36"><SPLITS/></RESULT><RESULT eventid="29" heatid="302" lane="7" points="327" resultid="2251" swimtime="00:02:43.98"><SPLITS><SPLIT distance="50" swimtime="00:00:34.43"/><SPLIT distance="100" swimtime="00:01:15.74"/><SPLIT distance="150" swimtime="00:01:59.66"/></SPLITS></RESULT><RESULT eventid="31" heatid="339" lane="5" points="290" resultid="2527" swimtime="00:01:36.85"><SPLITS><SPLIT distance="50" swimtime="00:00:45.37"/></SPLITS></RESULT><RESULT eventid="37" heatid="408" lane="7" points="338" resultid="3045" swimtime="00:02:57.01"><SPLITS><SPLIT distance="50" swimtime="00:00:41.67"/><SPLIT distance="100" swimtime="00:01:26.98"/><SPLIT distance="150" swimtime="00:02:13.63"/></SPLITS></RESULT><RESULT eventid="41" heatid="476" lane="4" points="323" resultid="3561" swimtime="00:06:27.99"><SPLITS><SPLIT distance="50" swimtime="00:00:42.30"/><SPLIT distance="100" swimtime="00:01:35.29"/><SPLIT distance="150" swimtime="00:02:24.36"/><SPLIT distance="200" swimtime="00:03:11.42"/><SPLIT distance="250" swimtime="00:04:06.00"/><SPLIT distance="300" swimtime="00:05:01.99"/><SPLIT distance="350" swimtime="00:05:45.74"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="267" birthdate="2010-01-01" firstname="Felix" gender="M" lastname="Adrion" license="411665"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="36" lane="1" points="207" resultid="267" swimtime="00:00:43.84"><SPLITS/></RESULT><RESULT eventid="6" heatid="74" lane="3" points="208" resultid="553" swimtime="00:01:23.36"><SPLITS><SPLIT distance="50" swimtime="00:00:36.75"/></SPLITS></RESULT><RESULT eventid="10" heatid="147" lane="8" points="286" resultid="1113" swimtime="00:00:31.72"><SPLITS/></RESULT><RESULT eventid="12" heatid="181" lane="7" points="242" resultid="1372" swimtime="00:03:02.76"><SPLITS><SPLIT distance="50" swimtime="00:00:36.51"/><SPLIT distance="100" swimtime="00:01:30.02"/><SPLIT distance="150" swimtime="00:02:23.08"/></SPLITS></RESULT><RESULT eventid="30" heatid="320" lane="8" points="274" resultid="2389" swimtime="00:02:36.90"><SPLITS><SPLIT distance="50" swimtime="00:00:33.97"/><SPLIT distance="100" swimtime="00:01:13.13"/><SPLIT distance="150" swimtime="00:01:55.85"/></SPLITS></RESULT><RESULT eventid="34" heatid="361" lane="7" points="171" resultid="2688" swimtime="00:03:18.78"><SPLITS><SPLIT distance="50" swimtime="00:00:38.01"/><SPLIT distance="100" swimtime="00:01:27.01"/><SPLIT distance="150" swimtime="00:02:21.82"/></SPLITS></RESULT><RESULT eventid="36" heatid="392" lane="5" points="233" resultid="2922" swimtime="00:00:36.17"><SPLITS/></RESULT><RESULT eventid="40" heatid="466" lane="2" points="275" resultid="3484" swimtime="00:01:12.03"><SPLITS><SPLIT distance="50" swimtime="00:00:33.77"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="274" birthdate="2011-01-01" firstname="Jonas" gender="M" lastname="Förtsch" license="435802"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="36" lane="8" points="236" resultid="274" swimtime="00:00:41.95"><SPLITS/></RESULT><RESULT eventid="8" heatid="97" lane="2" points="286" resultid="727" swimtime="00:03:11.02"><SPLITS><SPLIT distance="50" swimtime="00:00:43.81"/><SPLIT distance="100" swimtime="00:01:33.45"/><SPLIT distance="150" swimtime="00:02:22.59"/></SPLITS></RESULT><RESULT eventid="10" heatid="145" lane="8" points="224" resultid="1097" swimtime="00:00:34.43"><SPLITS/></RESULT><RESULT eventid="14" heatid="219" lane="7" points="190" resultid="1665" swimtime="00:01:29.72"><SPLITS><SPLIT distance="50" swimtime="00:00:43.24"/></SPLITS></RESULT><RESULT eventid="28" heatid="281" lane="1" points="194" resultid="2085" swimtime="00:00:40.90"><SPLITS/></RESULT><RESULT comment="12:52 Der Sportler führte mehr als den einen erlaubten kompletten Zyklus vollständig untergetaucht aus" eventid="32" heatid="352" lane="7" resultid="2625" status="DSQ" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="36" heatid="389" lane="3" points="167" resultid="2896" swimtime="00:00:40.40"><SPLITS/></RESULT><RESULT eventid="40" heatid="464" lane="3" points="247" resultid="3469" swimtime="00:01:14.59"><SPLITS><SPLIT distance="50" swimtime="00:00:36.59"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="279" birthdate="2007-01-01" firstname="Luca" gender="M" lastname="Schmidt" license="349907"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="37" lane="5" points="308" resultid="279" swimtime="00:00:38.42"><SPLITS/></RESULT><RESULT eventid="6" heatid="77" lane="7" points="344" resultid="581" swimtime="00:01:10.56"><SPLITS><SPLIT distance="50" swimtime="00:00:31.02"/></SPLITS></RESULT><RESULT eventid="10" heatid="152" lane="7" points="428" resultid="1152" swimtime="00:00:27.74"><SPLITS/></RESULT><RESULT eventid="14" heatid="223" lane="4" points="326" resultid="1693" swimtime="00:01:14.97"><SPLITS><SPLIT distance="50" swimtime="00:00:35.98"/></SPLITS></RESULT><RESULT eventid="28" heatid="286" lane="8" points="330" resultid="2131" swimtime="00:00:34.30"><SPLITS/></RESULT><RESULT eventid="32" heatid="354" lane="7" points="308" resultid="2641" swimtime="00:01:24.17"><SPLITS><SPLIT distance="50" swimtime="00:00:39.33"/></SPLITS></RESULT><RESULT eventid="36" heatid="395" lane="3" points="376" resultid="2944" swimtime="00:00:30.85"><SPLITS/></RESULT><RESULT eventid="40" heatid="470" lane="3" points="397" resultid="3516" swimtime="00:01:03.73"><SPLITS><SPLIT distance="50" swimtime="00:00:30.30"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="321" birthdate="2011-01-01" firstname="Lara" gender="F" lastname="Thelen" license="449401"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="43" lane="5" points="268" resultid="324" swimtime="00:06:06.52"><SPLITS><SPLIT distance="100" swimtime="00:01:27.92"/><SPLIT distance="200" swimtime="00:03:03.60"/><SPLIT distance="300" swimtime="00:04:37.31"/></SPLITS></RESULT><RESULT eventid="11" heatid="163" lane="3" points="272" resultid="1229" swimtime="00:03:14.55"><SPLITS><SPLIT distance="50" swimtime="00:00:45.45"/><SPLIT distance="100" swimtime="00:01:33.33"/><SPLIT distance="150" swimtime="00:02:31.96"/></SPLITS></RESULT><RESULT eventid="29" heatid="295" lane="4" points="283" resultid="2193" swimtime="00:02:51.94"><SPLITS><SPLIT distance="50" swimtime="00:00:38.38"/><SPLIT distance="100" swimtime="00:01:22.81"/><SPLIT distance="150" swimtime="00:02:08.55"/></SPLITS></RESULT><RESULT eventid="33" heatid="357" lane="4" points="188" resultid="2659" swimtime="00:03:32.28"><SPLITS><SPLIT distance="50" swimtime="00:00:44.71"/><SPLIT distance="100" swimtime="00:01:40.98"/><SPLIT distance="150" swimtime="00:02:37.69"/></SPLITS></RESULT><RESULT eventid="35" heatid="371" lane="7" points="208" resultid="2765" swimtime="00:00:41.18"><SPLITS/></RESULT><RESULT eventid="39" heatid="436" lane="1" points="277" resultid="3250" swimtime="00:01:19.29"><SPLITS><SPLIT distance="50" swimtime="00:00:38.79"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="344" birthdate="2011-01-01" firstname="Charlotte" gender="F" lastname="Karl" license="403795"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="48" lane="2" points="351" resultid="360" swimtime="00:05:35.03"><SPLITS><SPLIT distance="100" swimtime="00:01:17.06"/><SPLIT distance="200" swimtime="00:02:45.41"/><SPLIT distance="300" swimtime="00:04:12.29"/></SPLITS></RESULT><RESULT eventid="9" heatid="121" lane="4" points="386" resultid="915" swimtime="00:00:32.49"><SPLITS/></RESULT><RESULT eventid="13" heatid="205" lane="6" points="381" resultid="1557" swimtime="00:01:19.20"><SPLITS><SPLIT distance="50" swimtime="00:00:37.72"/></SPLITS></RESULT><RESULT eventid="27" heatid="270" lane="3" points="470" resultid="2005" swimtime="00:00:34.68"><SPLITS/></RESULT><RESULT eventid="31" heatid="338" lane="7" points="260" resultid="2521" swimtime="00:01:40.39"><SPLITS><SPLIT distance="50" swimtime="00:00:45.43"/></SPLITS></RESULT><RESULT eventid="37" heatid="410" lane="1" points="378" resultid="3055" swimtime="00:02:50.53"><SPLITS><SPLIT distance="50" swimtime="00:00:38.43"/><SPLIT distance="100" swimtime="00:01:21.85"/><SPLIT distance="150" swimtime="00:02:08.27"/></SPLITS></RESULT><RESULT eventid="39" heatid="443" lane="7" points="330" resultid="3311" swimtime="00:01:14.82"><SPLITS><SPLIT distance="50" swimtime="00:00:34.53"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="347" birthdate="2012-01-01" firstname="Valentina" gender="F" lastname="Ordnung" license="451809"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="48" lane="6" points="352" resultid="364" swimtime="00:05:34.72"><SPLITS><SPLIT distance="100" swimtime="00:01:18.72"/><SPLIT distance="200" swimtime="00:02:45.38"/><SPLIT distance="300" swimtime="00:04:13.22"/></SPLITS></RESULT><RESULT eventid="9" heatid="118" lane="6" points="360" resultid="893" swimtime="00:00:33.26"><SPLITS/></RESULT><RESULT eventid="13" heatid="200" lane="2" points="259" resultid="1513" swimtime="00:01:30.03"><SPLITS><SPLIT distance="50" swimtime="00:00:44.27"/></SPLITS></RESULT><RESULT eventid="29" heatid="300" lane="3" points="376" resultid="2232" swimtime="00:02:36.45"><SPLITS><SPLIT distance="50" swimtime="00:00:35.87"/><SPLIT distance="100" swimtime="00:01:15.14"/><SPLIT distance="150" swimtime="00:01:57.76"/></SPLITS></RESULT><RESULT eventid="35" heatid="370" lane="5" points="229" resultid="2755" swimtime="00:00:39.90"><SPLITS/></RESULT><RESULT eventid="39" heatid="439" lane="7" points="343" resultid="3280" swimtime="00:01:13.85"><SPLITS><SPLIT distance="50" swimtime="00:00:35.30"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="355" birthdate="2009-01-01" firstname="Dana" gender="F" lastname="Schörner" license="363135"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="49" lane="7" points="333" resultid="373" swimtime="00:05:40.98"><SPLITS><SPLIT distance="100" swimtime="00:01:14.61"/><SPLIT distance="200" swimtime="00:02:41.80"/><SPLIT distance="300" swimtime="00:04:12.11"/></SPLITS></RESULT><RESULT eventid="9" heatid="126" lane="5" points="458" resultid="956" swimtime="00:00:30.69"><SPLITS/></RESULT><RESULT eventid="13" heatid="202" lane="2" points="322" resultid="1529" swimtime="00:01:23.78"><SPLITS><SPLIT distance="50" swimtime="00:00:39.35"/></SPLITS></RESULT><RESULT eventid="27" heatid="268" lane="7" points="365" resultid="1994" swimtime="00:00:37.73"><SPLITS/></RESULT><RESULT eventid="29" heatid="303" lane="8" points="373" resultid="2260" swimtime="00:02:36.85"><SPLITS><SPLIT distance="50" swimtime="00:00:33.53"/><SPLIT distance="100" swimtime="00:01:12.05"/><SPLIT distance="150" swimtime="00:01:55.64"/></SPLITS></RESULT><RESULT eventid="35" heatid="378" lane="5" points="357" resultid="2816" swimtime="00:00:34.41"><SPLITS/></RESULT><RESULT eventid="39" heatid="445" lane="1" points="415" resultid="3321" swimtime="00:01:09.27"><SPLITS><SPLIT distance="50" swimtime="00:00:33.09"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="381" birthdate="2014-01-01" firstname="Ben" gender="M" lastname="Langheinrich" license="459878"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="54" lane="1" points="136" resultid="402" swimtime="00:07:07.00"><SPLITS><SPLIT distance="100" swimtime="00:01:36.06"/><SPLIT distance="200" swimtime="00:03:26.58"/><SPLIT distance="300" swimtime="00:05:21.25"/></SPLITS></RESULT><RESULT eventid="10" heatid="137" lane="8" points="120" resultid="1036" swimtime="00:00:42.30"><SPLITS/></RESULT><RESULT eventid="14" heatid="213" lane="2" points="131" resultid="1614" swimtime="00:01:41.48"><SPLITS><SPLIT distance="50" swimtime="00:00:50.55"/></SPLITS></RESULT><RESULT eventid="28" heatid="277" lane="5" points="110" resultid="2057" swimtime="00:00:49.47"><SPLITS/></RESULT><RESULT eventid="30" heatid="315" lane="1" points="130" resultid="2342" swimtime="00:03:21.13"><SPLITS><SPLIT distance="50" swimtime="00:00:45.20"/><SPLIT distance="100" swimtime="00:01:38.14"/><SPLIT distance="150" swimtime="00:02:32.09"/></SPLITS></RESULT><RESULT eventid="36" heatid="387" lane="3" points="53" resultid="2880" swimtime="00:00:59.06"><SPLITS/></RESULT><RESULT eventid="40" heatid="456" lane="1" points="112" resultid="3406" swimtime="00:01:37.05"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="388" birthdate="2013-01-01" firstname="Timur" gender="M" lastname="Gavlik" license="473447"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="55" lane="1" points="176" resultid="410" swimtime="00:06:32.29"><SPLITS><SPLIT distance="100" swimtime="00:01:25.93"/><SPLIT distance="200" swimtime="00:03:07.24"/><SPLIT distance="300" swimtime="00:04:51.67"/></SPLITS></RESULT><RESULT eventid="10" heatid="141" lane="7" points="163" resultid="1065" swimtime="00:00:38.26"><SPLITS/></RESULT><RESULT eventid="14" heatid="214" lane="2" points="137" resultid="1622" swimtime="00:01:40.08"><SPLITS><SPLIT distance="50" swimtime="00:00:48.17"/></SPLITS></RESULT><RESULT eventid="28" heatid="278" lane="2" points="148" resultid="2062" swimtime="00:00:44.77"><SPLITS/></RESULT><RESULT eventid="30" heatid="314" lane="6" points="170" resultid="2339" swimtime="00:03:04.03"><SPLITS><SPLIT distance="50" swimtime="00:00:38.18"/><SPLIT distance="100" swimtime="00:01:24.90"/><SPLIT distance="150" swimtime="00:02:15.90"/></SPLITS></RESULT><RESULT eventid="36" heatid="386" lane="7" points="74" resultid="2877" swimtime="00:00:52.83"><SPLITS/></RESULT><RESULT eventid="40" heatid="458" lane="3" points="164" resultid="3423" swimtime="00:01:25.57"><SPLITS><SPLIT distance="50" swimtime="00:00:41.72"/></SPLITS></RESULT></RESULTS></ATHLETE></ATHLETES><RELAYS/></CLUB><CLUB code="5085" name="SG Bamberg" nation="GER" region="02" shortname="Bamberg" type="CLUB"><CONTACT city="Bamberg" country="GER" email="coach@sgbamberg.de" name="Sikdar, Tushar" street="Steigerwaldstraße 9" zip="96049"/><OFFICIALS/><ATHLETES><ATHLETE athleteid="64" birthdate="2013-01-01" firstname="Emma" gender="F" lastname="Bauer" license="450240"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="9" lane="4" points="246" resultid="64" swimtime="00:00:46.74"><SPLITS/></RESULT><RESULT eventid="3" heatid="43" lane="7" points="227" resultid="326" swimtime="00:06:27.02"><SPLITS><SPLIT distance="100" swimtime="00:01:29.97"/><SPLIT distance="200" swimtime="00:03:10.90"/><SPLIT distance="300" swimtime="00:04:52.12"/></SPLITS></RESULT><RESULT eventid="11" heatid="163" lane="4" points="269" resultid="1230" swimtime="00:03:15.30"><SPLITS><SPLIT distance="50" swimtime="00:00:43.16"/><SPLIT distance="100" swimtime="00:01:33.83"/><SPLIT distance="150" swimtime="00:02:30.33"/></SPLITS></RESULT><RESULT eventid="13" heatid="198" lane="7" points="236" resultid="1502" swimtime="00:01:32.91"><SPLITS><SPLIT distance="50" swimtime="00:00:45.51"/></SPLITS></RESULT><RESULT eventid="19" heatid="235" lane="8" resultid="1769" swimtime="00:01:07.69"><SPLITS/></RESULT><RESULT eventid="29" heatid="295" lane="1" points="248" resultid="2190" swimtime="00:02:59.60"><SPLITS><SPLIT distance="50" swimtime="00:00:39.14"/><SPLIT distance="100" swimtime="00:01:24.24"/><SPLIT distance="150" swimtime="00:02:13.73"/></SPLITS></RESULT><RESULT eventid="37" heatid="405" lane="8" points="251" resultid="3022" swimtime="00:03:15.35"><SPLITS><SPLIT distance="50" swimtime="00:00:48.81"/><SPLIT distance="100" swimtime="00:01:38.59"/></SPLITS></RESULT><RESULT eventid="39" heatid="431" lane="3" points="262" resultid="3212" swimtime="00:01:20.80"><SPLITS><SPLIT distance="50" swimtime="00:00:38.71"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="68" birthdate="2014-01-01" firstname="Marie" gender="F" lastname="Glomb" license="450219"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="9" lane="8" points="226" resultid="68" swimtime="00:00:48.08"><SPLITS/></RESULT><RESULT eventid="3" heatid="42" lane="4" points="166" resultid="315" swimtime="00:07:09.29"><SPLITS><SPLIT distance="100" swimtime="00:01:35.44"/><SPLIT distance="200" swimtime="00:03:26.30"/><SPLIT distance="300" swimtime="00:05:18.89"/></SPLITS></RESULT><RESULT eventid="7" heatid="84" lane="2" points="229" resultid="626" swimtime="00:03:47.08"><SPLITS><SPLIT distance="50" swimtime="00:00:49.95"/><SPLIT distance="100" swimtime="00:01:46.93"/><SPLIT distance="150" swimtime="00:02:49.54"/></SPLITS></RESULT><RESULT eventid="11" heatid="159" lane="7" points="198" resultid="1201" swimtime="00:03:36.13"><SPLITS><SPLIT distance="50" swimtime="00:00:50.41"/><SPLIT distance="100" swimtime="00:01:49.89"/><SPLIT distance="150" swimtime="00:02:46.91"/></SPLITS></RESULT><RESULT eventid="25" heatid="248" lane="3" resultid="1839" swimtime="00:00:58.87"><SPLITS/></RESULT><RESULT eventid="31" heatid="335" lane="7" points="231" resultid="2497" swimtime="00:01:44.37"><SPLITS><SPLIT distance="50" swimtime="00:00:48.08"/></SPLITS></RESULT><RESULT eventid="35" heatid="365" lane="5" points="143" resultid="2715" swimtime="00:00:46.71"><SPLITS/></RESULT><RESULT eventid="39" heatid="428" lane="5" points="195" resultid="3190" swimtime="00:01:29.05"><SPLITS><SPLIT distance="50" swimtime="00:00:42.11"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="80" birthdate="2014-01-01" firstname="Lena" gender="F" lastname="Lempetzeder" license="450228"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="11" lane="4" resultid="80" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="3" heatid="43" lane="8" resultid="327" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="7" heatid="85" lane="5" resultid="637" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="11" heatid="159" lane="2" points="228" resultid="1197" swimtime="00:03:26.41"><SPLITS><SPLIT distance="50" swimtime="00:00:46.75"/><SPLIT distance="100" swimtime="00:01:38.04"/><SPLIT distance="150" swimtime="00:02:38.92"/></SPLITS></RESULT><RESULT eventid="25" heatid="248" lane="6" resultid="1842" swimtime="00:01:03.52"><SPLITS/></RESULT><RESULT eventid="31" heatid="333" lane="7" points="234" resultid="2481" swimtime="00:01:44.03"><SPLITS><SPLIT distance="50" swimtime="00:00:49.15"/></SPLITS></RESULT><RESULT eventid="35" heatid="366" lane="6" points="157" resultid="2724" swimtime="00:00:45.24"><SPLITS/></RESULT><RESULT eventid="39" heatid="428" lane="8" points="236" resultid="3193" swimtime="00:01:23.64"><SPLITS><SPLIT distance="50" swimtime="00:00:40.75"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="81" birthdate="2013-01-01" firstname="Katharina" gender="F" lastname="Dieter" license="446216"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="11" lane="5" points="253" resultid="81" swimtime="00:00:46.30"><SPLITS/></RESULT><RESULT eventid="3" heatid="42" lane="7" points="198" resultid="318" swimtime="00:06:45.15"><SPLITS><SPLIT distance="100" swimtime="00:01:29.22"/><SPLIT distance="200" swimtime="00:03:13.08"/><SPLIT distance="300" swimtime="00:05:00.55"/></SPLITS></RESULT><RESULT eventid="9" heatid="118" lane="3" points="359" resultid="890" swimtime="00:00:33.30"><SPLITS/></RESULT><RESULT eventid="11" heatid="162" lane="3" points="253" resultid="1221" swimtime="00:03:19.38"><SPLITS><SPLIT distance="50" swimtime="00:00:43.28"/><SPLIT distance="100" swimtime="00:01:37.90"/><SPLIT distance="150" swimtime="00:02:35.43"/></SPLITS></RESULT><RESULT eventid="23" heatid="242" lane="7" resultid="1805" swimtime="00:00:49.42"><SPLITS/></RESULT><RESULT eventid="29" heatid="295" lane="2" points="249" resultid="2191" swimtime="00:02:59.45"><SPLITS><SPLIT distance="50" swimtime="00:00:39.11"/><SPLIT distance="100" swimtime="00:01:24.12"/><SPLIT distance="150" swimtime="00:02:15.14"/></SPLITS></RESULT><RESULT eventid="35" heatid="368" lane="7" points="206" resultid="2741" swimtime="00:00:41.32"><SPLITS/></RESULT><RESULT eventid="39" heatid="433" lane="6" points="297" resultid="3231" swimtime="00:01:17.46"><SPLITS><SPLIT distance="50" swimtime="00:00:36.55"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="84" birthdate="2014-01-01" firstname="Hannah" gender="F" lastname="Bötsch" license="461183"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="11" lane="8" points="196" resultid="84" swimtime="00:00:50.38"><SPLITS/></RESULT><RESULT eventid="3" heatid="45" lane="1" points="298" resultid="336" swimtime="00:05:53.90"><SPLITS><SPLIT distance="100" swimtime="00:01:22.06"/><SPLIT distance="200" swimtime="00:02:52.58"/><SPLIT distance="300" swimtime="00:04:24.75"/></SPLITS></RESULT><RESULT eventid="11" heatid="165" lane="2" points="282" resultid="1244" swimtime="00:03:12.11"><SPLITS><SPLIT distance="50" swimtime="00:00:42.82"/><SPLIT distance="100" swimtime="00:01:31.68"/><SPLIT distance="150" swimtime="00:02:30.81"/></SPLITS></RESULT><RESULT eventid="13" heatid="198" lane="2" points="215" resultid="1497" swimtime="00:01:35.81"><SPLITS><SPLIT distance="50" swimtime="00:00:48.55"/></SPLITS></RESULT><RESULT eventid="23" heatid="243" lane="8" resultid="1814" swimtime="00:00:50.26"><SPLITS/></RESULT><RESULT eventid="29" heatid="297" lane="4" points="322" resultid="2209" swimtime="00:02:44.68"><SPLITS><SPLIT distance="50" swimtime="00:00:37.74"/><SPLIT distance="100" swimtime="00:01:20.72"/><SPLIT distance="150" swimtime="00:02:03.62"/></SPLITS></RESULT><RESULT eventid="35" heatid="369" lane="3" points="228" resultid="2745" swimtime="00:00:39.96"><SPLITS/></RESULT><RESULT eventid="39" heatid="434" lane="3" points="294" resultid="3236" swimtime="00:01:17.69"><SPLITS><SPLIT distance="50" swimtime="00:00:38.40"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="109" birthdate="2010-01-01" firstname="Hannah" gender="F" lastname="Drescher" license="410251"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="15" lane="1" points="234" resultid="109" swimtime="00:00:47.53"><SPLITS/></RESULT><RESULT eventid="3" heatid="47" lane="7" points="318" resultid="358" swimtime="00:05:46.03"><SPLITS><SPLIT distance="100" swimtime="00:01:17.84"/><SPLIT distance="200" swimtime="00:02:47.27"/><SPLIT distance="300" swimtime="00:04:18.40"/></SPLITS></RESULT><RESULT eventid="9" heatid="119" lane="2" points="330" resultid="897" swimtime="00:00:34.22"><SPLITS/></RESULT><RESULT eventid="11" heatid="166" lane="8" points="294" resultid="1258" swimtime="00:03:09.56"><SPLITS><SPLIT distance="50" swimtime="00:00:42.97"/><SPLIT distance="100" swimtime="00:01:28.53"/><SPLIT distance="150" swimtime="00:02:28.37"/></SPLITS></RESULT><RESULT eventid="27" heatid="262" lane="1" points="294" resultid="1940" swimtime="00:00:40.57"><SPLITS/></RESULT><RESULT eventid="29" heatid="300" lane="7" points="343" resultid="2236" swimtime="00:02:41.36"><SPLITS><SPLIT distance="50" swimtime="00:00:36.16"/><SPLIT distance="100" swimtime="00:01:17.48"/><SPLIT distance="150" swimtime="00:01:59.93"/></SPLITS></RESULT><RESULT eventid="35" heatid="369" lane="6" points="197" resultid="2748" swimtime="00:00:41.97"><SPLITS/></RESULT><RESULT eventid="39" heatid="438" lane="8" points="311" resultid="3273" swimtime="00:01:16.26"><SPLITS><SPLIT distance="50" swimtime="00:00:37.19"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="122" birthdate="2011-01-01" firstname="Emily" gender="F" lastname="Liedtke" license="441612"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="16" lane="6" points="317" resultid="122" swimtime="00:00:42.95"><SPLITS/></RESULT><RESULT eventid="3" heatid="49" lane="6" points="398" resultid="372" swimtime="00:05:21.20"><SPLITS><SPLIT distance="100" swimtime="00:01:14.99"/><SPLIT distance="200" swimtime="00:02:40.95"/><SPLIT distance="300" swimtime="00:04:05.70"/></SPLITS></RESULT><RESULT eventid="9" heatid="125" lane="7" points="435" resultid="950" swimtime="00:00:31.22"><SPLITS/></RESULT><RESULT eventid="11" heatid="168" lane="6" points="366" resultid="1272" swimtime="00:02:56.18"><SPLITS><SPLIT distance="50" swimtime="00:00:39.73"/><SPLIT distance="100" swimtime="00:01:25.46"/><SPLIT distance="150" swimtime="00:02:19.07"/></SPLITS></RESULT><RESULT eventid="27" heatid="262" lane="6" points="376" resultid="1945" swimtime="00:00:37.36"><SPLITS/></RESULT><RESULT eventid="29" heatid="301" lane="2" points="452" resultid="2239" swimtime="00:02:27.16"><SPLITS><SPLIT distance="50" swimtime="00:00:33.93"/><SPLIT distance="100" swimtime="00:01:13.05"/><SPLIT distance="150" swimtime="00:01:51.67"/></SPLITS></RESULT><RESULT eventid="35" heatid="372" lane="6" points="265" resultid="2772" swimtime="00:00:37.99"><SPLITS/></RESULT><RESULT eventid="39" heatid="442" lane="2" points="452" resultid="3298" swimtime="00:01:07.34"><SPLITS><SPLIT distance="50" swimtime="00:00:32.28"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="124" birthdate="2014-01-01" firstname="Hailey" gender="F" lastname="Heron" license="474925"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="16" lane="8" points="197" resultid="124" swimtime="00:00:50.29"><SPLITS/></RESULT><RESULT eventid="3" heatid="44" lane="3" points="260" resultid="330" swimtime="00:06:10.20"><SPLITS><SPLIT distance="100" swimtime="00:01:26.41"/><SPLIT distance="200" swimtime="00:03:02.16"/><SPLIT distance="300" swimtime="00:04:37.70"/></SPLITS></RESULT><RESULT eventid="9" heatid="118" lane="7" points="321" resultid="894" swimtime="00:00:34.55"><SPLITS/></RESULT><RESULT eventid="11" heatid="164" lane="2" resultid="1236" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="23" heatid="242" lane="4" resultid="1802" swimtime="00:00:51.70"><SPLITS/></RESULT><RESULT eventid="29" heatid="297" lane="5" points="294" resultid="2210" swimtime="00:02:49.89"><SPLITS><SPLIT distance="50" swimtime="00:00:38.75"/><SPLIT distance="100" swimtime="00:01:22.72"/><SPLIT distance="150" swimtime="00:02:07.43"/></SPLITS></RESULT><RESULT eventid="35" heatid="371" lane="8" points="227" resultid="2766" swimtime="00:00:40.04"><SPLITS/></RESULT><RESULT eventid="39" heatid="436" lane="6" points="323" resultid="3255" swimtime="00:01:15.31"><SPLITS><SPLIT distance="50" swimtime="00:00:35.54"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="129" birthdate="2009-01-01" firstname="Olivia" gender="F" lastname="Lange" license="398680"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="17" lane="5" resultid="129" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="5" heatid="69" lane="2" resultid="513" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="9" heatid="124" lane="3" resultid="938" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="27" heatid="266" lane="4" resultid="1975" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="35" heatid="379" lane="8" resultid="2827" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="39" heatid="445" lane="7" resultid="3327" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="138" birthdate="2011-01-01" firstname="Eva" gender="F" lastname="Jakubaß" license="409223"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="18" lane="6" points="290" resultid="138" swimtime="00:00:44.24"><SPLITS/></RESULT><RESULT eventid="3" heatid="50" lane="3" points="406" resultid="377" swimtime="00:05:19.15"><SPLITS><SPLIT distance="100" swimtime="00:01:15.00"/><SPLIT distance="200" swimtime="00:02:36.25"/><SPLIT distance="300" swimtime="00:03:58.62"/></SPLITS></RESULT><RESULT eventid="9" heatid="125" lane="8" points="398" resultid="951" swimtime="00:00:32.16"><SPLITS/></RESULT><RESULT eventid="17" heatid="231" lane="3" points="415" resultid="1742" swimtime="00:10:49.92"><SPLITS><SPLIT distance="100" swimtime="00:01:15.04"/><SPLIT distance="200" swimtime="00:02:36.67"/><SPLIT distance="300" swimtime="00:03:58.47"/><SPLIT distance="400" swimtime="00:05:21.58"/><SPLIT distance="500" swimtime="00:06:44.28"/><SPLIT distance="600" swimtime="00:08:07.66"/><SPLIT distance="700" swimtime="00:09:30.08"/></SPLITS></RESULT><RESULT eventid="31" heatid="340" lane="1" points="286" resultid="2531" swimtime="00:01:37.27"><SPLITS><SPLIT distance="50" swimtime="00:00:46.37"/></SPLITS></RESULT><RESULT eventid="39" heatid="446" lane="4" points="426" resultid="3331" swimtime="00:01:08.70"><SPLITS><SPLIT distance="50" swimtime="00:00:32.30"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="155" birthdate="2011-01-01" firstname="Eva" gender="F" lastname="Meister" license="409222"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="20" lane="7" points="387" resultid="155" swimtime="00:00:40.18"><SPLITS/></RESULT><RESULT eventid="9" heatid="120" lane="7" points="432" resultid="910" swimtime="00:00:31.29"><SPLITS/></RESULT><RESULT eventid="17" heatid="230" lane="4" points="341" resultid="1735" swimtime="00:11:33.72"><SPLITS><SPLIT distance="100" swimtime="00:01:19.53"/><SPLIT distance="200" swimtime="00:02:47.40"/><SPLIT distance="300" swimtime="00:04:16.05"/><SPLIT distance="400" swimtime="00:05:46.18"/><SPLIT distance="500" swimtime="00:07:15.33"/><SPLIT distance="600" swimtime="00:08:43.98"/><SPLIT distance="700" swimtime="00:10:11.69"/></SPLITS></RESULT><RESULT eventid="31" heatid="340" lane="4" points="362" resultid="2534" swimtime="00:01:29.96"><SPLITS><SPLIT distance="50" swimtime="00:00:40.61"/></SPLITS></RESULT><RESULT eventid="35" heatid="374" lane="4" points="365" resultid="2786" swimtime="00:00:34.17"><SPLITS/></RESULT><RESULT eventid="39" heatid="441" lane="7" points="398" resultid="3295" swimtime="00:01:10.29"><SPLITS><SPLIT distance="50" swimtime="00:00:32.84"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="160" birthdate="2011-01-01" firstname="Mara" gender="F" lastname="Friedemann" license="434413"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="21" lane="4" points="416" resultid="160" swimtime="00:00:39.24"><SPLITS/></RESULT><RESULT eventid="7" heatid="89" lane="7" points="325" resultid="671" swimtime="00:03:22.02"><SPLITS><SPLIT distance="50" swimtime="00:00:45.16"/><SPLIT distance="100" swimtime="00:01:37.63"/><SPLIT distance="150" swimtime="00:02:29.51"/></SPLITS></RESULT><RESULT eventid="9" heatid="127" lane="8" points="415" resultid="966" swimtime="00:00:31.71"><SPLITS/></RESULT><RESULT eventid="29" heatid="302" lane="1" points="382" resultid="2245" swimtime="00:02:35.63"><SPLITS><SPLIT distance="50" swimtime="00:00:34.03"/><SPLIT distance="100" swimtime="00:01:13.33"/><SPLIT distance="150" swimtime="00:01:55.64"/></SPLITS></RESULT><RESULT eventid="31" heatid="341" lane="8" points="337" resultid="2546" swimtime="00:01:32.09"><SPLITS><SPLIT distance="50" swimtime="00:00:43.12"/></SPLITS></RESULT><RESULT eventid="39" heatid="444" lane="7" points="405" resultid="3319" swimtime="00:01:09.87"><SPLITS><SPLIT distance="50" swimtime="00:00:32.99"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="221" birthdate="2013-01-01" firstname="Ferdinand" gender="M" lastname="Krome" license="446214"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="30" lane="1" points="136" resultid="221" swimtime="00:00:50.41"><SPLITS/></RESULT><RESULT eventid="4" heatid="56" lane="5" points="204" resultid="422" swimtime="00:06:13.83"><SPLITS><SPLIT distance="100" swimtime="00:01:26.25"/><SPLIT distance="200" swimtime="00:03:02.30"/><SPLIT distance="300" swimtime="00:04:38.79"/></SPLITS></RESULT><RESULT eventid="12" heatid="178" lane="3" points="166" resultid="1344" swimtime="00:03:27.15"><SPLITS><SPLIT distance="50" swimtime="00:00:50.70"/><SPLIT distance="100" swimtime="00:01:41.88"/><SPLIT distance="150" swimtime="00:02:44.57"/></SPLITS></RESULT><RESULT eventid="14" heatid="215" lane="8" points="158" resultid="1634" swimtime="00:01:35.30"><SPLITS><SPLIT distance="50" swimtime="00:00:48.69"/></SPLITS></RESULT><RESULT eventid="24" heatid="245" lane="7" resultid="1826" swimtime="00:00:57.54"><SPLITS/></RESULT><RESULT eventid="30" heatid="315" lane="3" points="194" resultid="2344" swimtime="00:02:55.92"><SPLITS><SPLIT distance="50" swimtime="00:00:39.43"/><SPLIT distance="100" swimtime="00:01:24.16"/><SPLIT distance="150" swimtime="00:02:11.30"/></SPLITS></RESULT><RESULT eventid="36" heatid="386" lane="3" points="110" resultid="2873" swimtime="00:00:46.36"><SPLITS/></RESULT><RESULT eventid="40" heatid="460" lane="8" points="183" resultid="3443" swimtime="00:01:22.41"><SPLITS><SPLIT distance="50" swimtime="00:00:39.20"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="252" birthdate="2013-01-01" firstname="Thomas" gender="M" lastname="Kraus" license="456925"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="33" lane="8" points="171" resultid="252" swimtime="00:00:46.68"><SPLITS/></RESULT><RESULT eventid="4" heatid="56" lane="4" points="212" resultid="421" swimtime="00:06:08.64"><SPLITS><SPLIT distance="100" swimtime="00:01:25.94"/><SPLIT distance="200" swimtime="00:03:02.26"/><SPLIT distance="300" swimtime="00:04:38.13"/></SPLITS></RESULT><RESULT eventid="10" heatid="144" lane="5" points="234" resultid="1086" swimtime="00:00:33.90"><SPLITS/></RESULT><RESULT eventid="12" heatid="178" lane="4" points="176" resultid="1345" swimtime="00:03:23.42"><SPLITS><SPLIT distance="50" swimtime="00:00:47.76"/><SPLIT distance="100" swimtime="00:01:44.52"/><SPLIT distance="150" swimtime="00:02:42.31"/></SPLITS></RESULT><RESULT eventid="24" heatid="245" lane="8" resultid="1827" swimtime="00:00:56.41"><SPLITS/></RESULT><RESULT eventid="30" heatid="315" lane="4" points="208" resultid="2345" swimtime="00:02:52.00"><SPLITS><SPLIT distance="50" swimtime="00:00:37.88"/><SPLIT distance="100" swimtime="00:01:23.54"/><SPLIT distance="150" swimtime="00:02:09.41"/></SPLITS></RESULT><RESULT eventid="36" heatid="385" lane="4" points="144" resultid="2866" swimtime="00:00:42.47"><SPLITS/></RESULT><RESULT eventid="40" heatid="463" lane="2" points="245" resultid="3461" swimtime="00:01:14.88"><SPLITS><SPLIT distance="50" swimtime="00:00:35.43"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="258" birthdate="2011-01-01" firstname="Christopher" gender="M" lastname="Flach" license="443319"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="34" lane="6" points="235" resultid="258" swimtime="00:00:42.01"><SPLITS/></RESULT><RESULT eventid="4" heatid="58" lane="1" points="233" resultid="434" swimtime="00:05:57.16"><SPLITS><SPLIT distance="100" swimtime="00:01:18.56"/><SPLIT distance="200" swimtime="00:02:50.41"/><SPLIT distance="300" swimtime="00:04:24.56"/></SPLITS></RESULT><RESULT eventid="12" heatid="181" lane="8" points="226" resultid="1373" swimtime="00:03:06.91"><SPLITS><SPLIT distance="50" swimtime="00:00:43.51"/><SPLIT distance="100" swimtime="00:01:30.51"/><SPLIT distance="150" swimtime="00:02:25.33"/></SPLITS></RESULT><RESULT eventid="14" heatid="219" lane="2" points="190" resultid="1660" swimtime="00:01:29.60"><SPLITS><SPLIT distance="50" swimtime="00:00:43.13"/></SPLITS></RESULT><RESULT eventid="28" heatid="281" lane="2" points="192" resultid="2086" swimtime="00:00:41.07"><SPLITS/></RESULT><RESULT eventid="30" heatid="317" lane="4" points="225" resultid="2361" swimtime="00:02:47.59"><SPLITS><SPLIT distance="50" swimtime="00:00:35.53"/><SPLIT distance="100" swimtime="00:01:18.40"/><SPLIT distance="150" swimtime="00:02:03.35"/></SPLITS></RESULT><RESULT eventid="38" heatid="416" lane="7" points="204" resultid="3105" swimtime="00:03:10.03"><SPLITS><SPLIT distance="50" swimtime="00:00:43.07"/><SPLIT distance="100" swimtime="00:01:31.66"/><SPLIT distance="150" swimtime="00:02:21.55"/></SPLITS></RESULT><RESULT eventid="40" heatid="462" lane="2" points="211" resultid="3453" swimtime="00:01:18.61"><SPLITS><SPLIT distance="50" swimtime="00:00:36.64"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="262" birthdate="2009-01-01" firstname="Robert" gender="M" lastname="Hartmann" license="377373"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="35" lane="4" points="422" resultid="262" swimtime="00:00:34.57"><SPLITS/></RESULT><RESULT eventid="10" heatid="155" lane="3" points="529" resultid="1171" swimtime="00:00:25.85"><SPLITS/></RESULT><RESULT eventid="12" heatid="188" lane="7" points="473" resultid="1426" swimtime="00:02:26.23"><SPLITS><SPLIT distance="50" swimtime="00:00:30.43"/><SPLIT distance="100" swimtime="00:01:09.32"/><SPLIT distance="150" swimtime="00:01:54.33"/></SPLITS></RESULT><RESULT eventid="28" heatid="286" lane="4" points="497" resultid="2127" swimtime="00:00:29.93"><SPLITS/></RESULT><RESULT eventid="36" heatid="398" lane="7" points="522" resultid="2972" swimtime="00:00:27.65"><SPLITS/></RESULT><RESULT eventid="40" heatid="474" lane="2" points="607" resultid="3546" swimtime="00:00:55.34"><SPLITS><SPLIT distance="50" swimtime="00:00:26.45"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="276" birthdate="2009-01-01" firstname="Raphael" gender="M" lastname="Jakubaß" license="392827"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="37" lane="2" points="347" resultid="276" swimtime="00:00:36.90"><SPLITS/></RESULT><RESULT eventid="8" heatid="100" lane="7" points="375" resultid="755" swimtime="00:02:54.56"><SPLITS><SPLIT distance="50" swimtime="00:00:38.89"/><SPLIT distance="100" swimtime="00:01:24.11"/><SPLIT distance="150" swimtime="00:02:08.00"/></SPLITS></RESULT><RESULT eventid="12" heatid="186" lane="5" points="379" resultid="1408" swimtime="00:02:37.46"><SPLITS><SPLIT distance="50" swimtime="00:00:33.46"/><SPLIT distance="100" swimtime="00:01:16.70"/><SPLIT distance="150" swimtime="00:02:01.28"/></SPLITS></RESULT><RESULT eventid="30" heatid="322" lane="6" points="409" resultid="2401" swimtime="00:02:17.41"><SPLITS><SPLIT distance="50" swimtime="00:00:31.34"/><SPLIT distance="100" swimtime="00:01:05.80"/><SPLIT distance="150" swimtime="00:01:42.07"/></SPLITS></RESULT><RESULT eventid="32" heatid="353" lane="4" points="366" resultid="2630" swimtime="00:01:19.45"><SPLITS><SPLIT distance="50" swimtime="00:00:36.88"/></SPLITS></RESULT><RESULT eventid="40" heatid="469" lane="8" points="413" resultid="3513" swimtime="00:01:02.89"><SPLITS><SPLIT distance="50" swimtime="00:00:31.01"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="282" birthdate="2011-01-01" firstname="Raphael" gender="M" lastname="Erhard" license="477014"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="37" lane="8" points="401" resultid="282" swimtime="00:00:35.18"><SPLITS/></RESULT><RESULT eventid="6" heatid="76" lane="8" points="374" resultid="574" swimtime="00:01:08.59"><SPLITS><SPLIT distance="50" swimtime="00:00:32.13"/></SPLITS></RESULT><RESULT eventid="10" heatid="153" lane="2" points="495" resultid="1155" swimtime="00:00:26.42"><SPLITS/></RESULT><RESULT eventid="12" heatid="187" lane="2" points="438" resultid="1413" swimtime="00:02:30.03"><SPLITS><SPLIT distance="50" swimtime="00:00:31.28"/><SPLIT distance="100" swimtime="00:01:10.81"/><SPLIT distance="150" swimtime="00:01:57.01"/></SPLITS></RESULT><RESULT eventid="32" heatid="353" lane="6" points="412" resultid="2632" swimtime="00:01:16.42"><SPLITS><SPLIT distance="50" swimtime="00:00:36.36"/></SPLITS></RESULT><RESULT eventid="36" heatid="393" lane="6" points="471" resultid="2931" swimtime="00:00:28.61"><SPLITS/></RESULT><RESULT eventid="40" heatid="473" lane="7" points="540" resultid="3543" swimtime="00:00:57.52"><SPLITS><SPLIT distance="50" swimtime="00:00:28.21"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="297" birthdate="2010-01-01" firstname="Szymon" gender="M" lastname="Gorczynski" license="409225"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="39" lane="7" points="472" resultid="297" swimtime="00:00:33.32"><SPLITS/></RESULT><RESULT eventid="8" heatid="100" lane="6" points="425" resultid="754" swimtime="00:02:47.40"><SPLITS><SPLIT distance="50" swimtime="00:00:37.49"/><SPLIT distance="100" swimtime="00:01:20.92"/><SPLIT distance="150" swimtime="00:02:02.79"/></SPLITS></RESULT><RESULT eventid="10" heatid="149" lane="6" points="372" resultid="1127" swimtime="00:00:29.07"><SPLITS/></RESULT><RESULT eventid="32" heatid="355" lane="7" points="417" resultid="2648" swimtime="00:01:16.12"><SPLITS><SPLIT distance="50" swimtime="00:00:34.77"/></SPLITS></RESULT><RESULT eventid="36" heatid="394" lane="7" points="294" resultid="2940" swimtime="00:00:33.47"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="312" birthdate="2013-01-01" firstname="Anni" gender="F" lastname="Kreis" license="450215"><HANDICAP/><ENTRIES/><RESULTS><RESULT comment="10:09 Die Schwimmerin hat wiederholt die Startbahn gewechselt" eventid="3" heatid="42" lane="2" resultid="313" status="DSQ" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="5" heatid="63" lane="6" points="178" resultid="472" swimtime="00:01:38.61"><SPLITS><SPLIT distance="50" swimtime="00:00:45.96"/></SPLITS></RESULT><RESULT eventid="11" heatid="162" lane="5" points="272" resultid="1223" swimtime="00:03:14.65"><SPLITS><SPLIT distance="50" swimtime="00:00:44.42"/><SPLIT distance="100" swimtime="00:01:32.50"/><SPLIT distance="150" swimtime="00:02:31.27"/></SPLITS></RESULT><RESULT eventid="13" heatid="197" lane="3" points="231" resultid="1490" swimtime="00:01:33.63"><SPLITS><SPLIT distance="50" swimtime="00:00:46.98"/></SPLITS></RESULT><RESULT eventid="23" heatid="242" lane="1" resultid="1799" swimtime="00:00:53.56"><SPLITS/></RESULT><RESULT eventid="29" heatid="294" lane="6" points="240" resultid="2187" swimtime="00:03:01.58"><SPLITS><SPLIT distance="50" swimtime="00:00:40.04"/><SPLIT distance="100" swimtime="00:01:27.58"/><SPLIT distance="150" swimtime="00:02:16.23"/></SPLITS></RESULT><RESULT eventid="35" heatid="370" lane="7" points="230" resultid="2757" swimtime="00:00:39.82"><SPLITS/></RESULT><RESULT eventid="39" heatid="433" lane="7" points="259" resultid="3232" swimtime="00:01:21.10"><SPLITS><SPLIT distance="50" swimtime="00:00:37.46"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="314" birthdate="2013-01-01" firstname="Ella" gender="F" lastname="Schaubert" license="446457"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="42" lane="5" resultid="316" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="7" heatid="87" lane="8" resultid="656" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="11" heatid="162" lane="7" resultid="1225" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="13" heatid="196" lane="5" points="149" resultid="1484" swimtime="00:01:48.31"><SPLITS/></RESULT><RESULT eventid="25" heatid="248" lane="2" resultid="1838" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="31" heatid="336" lane="1" resultid="2499" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="35" heatid="370" lane="3" resultid="2753" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="39" heatid="432" lane="7" resultid="3224" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="317" birthdate="2012-01-01" firstname="Bella Victoria" gender="F" lastname="Kostylieva" license="437501"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="43" lane="1" points="226" resultid="320" swimtime="00:06:27.65"><SPLITS><SPLIT distance="100" swimtime="00:01:27.49"/><SPLIT distance="200" swimtime="00:03:09.00"/><SPLIT distance="300" swimtime="00:04:51.15"/></SPLITS></RESULT><RESULT eventid="5" heatid="64" lane="2" points="116" resultid="474" swimtime="00:01:53.57"><SPLITS><SPLIT distance="50" swimtime="00:00:49.43"/></SPLITS></RESULT><RESULT eventid="9" heatid="113" lane="2" points="242" resultid="850" swimtime="00:00:37.97"><SPLITS/></RESULT><RESULT eventid="11" heatid="161" lane="3" points="234" resultid="1213" swimtime="00:03:24.47"><SPLITS><SPLIT distance="50" swimtime="00:00:50.68"/><SPLIT distance="100" swimtime="00:01:45.24"/><SPLIT distance="150" swimtime="00:02:40.93"/></SPLITS></RESULT><RESULT eventid="27" heatid="258" lane="4" points="255" resultid="1911" swimtime="00:00:42.54"><SPLITS/></RESULT><RESULT eventid="29" heatid="294" lane="4" points="218" resultid="2185" swimtime="00:03:07.44"><SPLITS><SPLIT distance="50" swimtime="00:00:40.46"/><SPLIT distance="100" swimtime="00:01:29.30"/><SPLIT distance="150" swimtime="00:02:18.89"/></SPLITS></RESULT><RESULT eventid="37" heatid="404" lane="8" points="234" resultid="3014" swimtime="00:03:20.03"><SPLITS><SPLIT distance="50" swimtime="00:00:49.02"/><SPLIT distance="100" swimtime="00:01:40.61"/><SPLIT distance="150" swimtime="00:02:33.52"/></SPLITS></RESULT><RESULT eventid="39" heatid="430" lane="4" points="240" resultid="3205" swimtime="00:01:23.16"><SPLITS><SPLIT distance="50" swimtime="00:00:38.92"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="320" birthdate="2014-01-01" firstname="Charlotte" gender="F" lastname="Müller-Bergh" license="468708"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="43" lane="4" points="235" resultid="323" swimtime="00:06:22.66"><SPLITS><SPLIT distance="100" swimtime="00:01:28.56"/><SPLIT distance="200" swimtime="00:03:07.48"/><SPLIT distance="300" swimtime="00:04:47.76"/></SPLITS></RESULT><RESULT eventid="7" heatid="88" lane="3" points="243" resultid="659" swimtime="00:03:42.55"><SPLITS><SPLIT distance="50" swimtime="00:00:52.64"/><SPLIT distance="100" swimtime="00:01:47.71"/><SPLIT distance="150" swimtime="00:02:47.01"/></SPLITS></RESULT><RESULT eventid="11" heatid="164" lane="4" resultid="1238" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="13" heatid="195" lane="5" resultid="1476" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="25" heatid="249" lane="3" resultid="1847" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="31" heatid="338" lane="8" resultid="2522" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="37" heatid="403" lane="1" resultid="2999" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="39" heatid="432" lane="4" resultid="3221" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="323" birthdate="2011-01-01" firstname="Lara" gender="F" lastname="Hünniger" license="425312"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="44" lane="1" points="282" resultid="328" swimtime="00:06:00.28"><SPLITS><SPLIT distance="100" swimtime="00:01:20.65"/><SPLIT distance="200" swimtime="00:02:51.94"/><SPLIT distance="300" swimtime="00:04:26.00"/></SPLITS></RESULT><RESULT eventid="7" heatid="87" lane="6" points="320" resultid="654" swimtime="00:03:22.97"><SPLITS><SPLIT distance="50" swimtime="00:00:44.31"/><SPLIT distance="100" swimtime="00:01:35.03"/><SPLIT distance="150" swimtime="00:02:28.98"/></SPLITS></RESULT><RESULT eventid="11" heatid="163" lane="5" points="318" resultid="1231" swimtime="00:03:04.71"><SPLITS><SPLIT distance="50" swimtime="00:00:42.37"/><SPLIT distance="100" swimtime="00:01:30.75"/><SPLIT distance="150" swimtime="00:02:23.86"/></SPLITS></RESULT><RESULT eventid="29" heatid="296" lane="1" points="340" resultid="2198" swimtime="00:02:41.83"><SPLITS><SPLIT distance="50" swimtime="00:00:37.45"/><SPLIT distance="100" swimtime="00:01:18.84"/><SPLIT distance="150" swimtime="00:02:02.92"/></SPLITS></RESULT><RESULT eventid="31" heatid="340" lane="8" points="340" resultid="2538" swimtime="00:01:31.85"><SPLITS><SPLIT distance="50" swimtime="00:00:45.07"/></SPLITS></RESULT><RESULT eventid="35" heatid="370" lane="1" points="252" resultid="2751" swimtime="00:00:38.67"><SPLITS/></RESULT><RESULT eventid="39" heatid="434" lane="5" points="393" resultid="3238" swimtime="00:01:10.59"><SPLITS><SPLIT distance="50" swimtime="00:00:35.00"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="324" birthdate="2010-01-01" firstname="Alina" gender="F" lastname="Lotar" license="406867"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="44" lane="2" points="309" resultid="329" swimtime="00:05:49.48"><SPLITS><SPLIT distance="100" swimtime="00:01:21.29"/><SPLIT distance="200" swimtime="00:02:51.37"/><SPLIT distance="300" swimtime="00:04:22.49"/></SPLITS></RESULT><RESULT eventid="5" heatid="65" lane="1" points="212" resultid="481" swimtime="00:01:32.95"><SPLITS><SPLIT distance="50" swimtime="00:00:41.26"/></SPLITS></RESULT><RESULT eventid="9" heatid="117" lane="6" points="319" resultid="885" swimtime="00:00:34.62"><SPLITS/></RESULT><RESULT eventid="11" heatid="165" lane="6" points="313" resultid="1248" swimtime="00:03:05.65"><SPLITS><SPLIT distance="50" swimtime="00:00:40.86"/><SPLIT distance="100" swimtime="00:01:29.52"/><SPLIT distance="150" swimtime="00:02:22.69"/></SPLITS></RESULT><RESULT eventid="33" heatid="357" lane="3" points="185" resultid="2658" swimtime="00:03:33.73"><SPLITS><SPLIT distance="50" swimtime="00:00:43.12"/><SPLIT distance="100" swimtime="00:01:36.41"/><SPLIT distance="150" swimtime="00:02:35.99"/></SPLITS></RESULT><RESULT eventid="35" heatid="370" lane="8" points="210" resultid="2758" swimtime="00:00:41.04"><SPLITS/></RESULT><RESULT eventid="39" heatid="435" lane="7" points="309" resultid="3248" swimtime="00:01:16.41"><SPLITS><SPLIT distance="50" swimtime="00:00:36.73"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="334" birthdate="2012-01-01" firstname="Lena" gender="F" lastname="Troll" license="438002"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="45" lane="7" points="315" resultid="342" swimtime="00:05:47.17"><SPLITS><SPLIT distance="200" swimtime="00:02:50.21"/><SPLIT distance="300" swimtime="00:04:20.12"/></SPLITS></RESULT><RESULT eventid="7" heatid="87" lane="1" points="335" resultid="649" swimtime="00:03:19.97"><SPLITS><SPLIT distance="50" swimtime="00:00:45.50"/><SPLIT distance="100" swimtime="00:01:35.79"/><SPLIT distance="150" swimtime="00:02:30.60"/></SPLITS></RESULT><RESULT eventid="9" heatid="124" lane="8" points="403" resultid="943" swimtime="00:00:32.02"><SPLITS/></RESULT><RESULT eventid="11" heatid="167" lane="4" points="347" resultid="1262" swimtime="00:02:59.33"><SPLITS><SPLIT distance="50" swimtime="00:00:40.96"/><SPLIT distance="100" swimtime="00:01:27.88"/><SPLIT distance="150" swimtime="00:02:19.16"/></SPLITS></RESULT><RESULT eventid="29" heatid="298" lane="8" points="354" resultid="2221" swimtime="00:02:39.61"><SPLITS><SPLIT distance="50" swimtime="00:00:38.31"/><SPLIT distance="100" swimtime="00:01:18.42"/><SPLIT distance="150" swimtime="00:02:01.16"/></SPLITS></RESULT><RESULT eventid="31" heatid="339" lane="4" points="326" resultid="2526" swimtime="00:01:33.15"><SPLITS><SPLIT distance="50" swimtime="00:00:43.42"/></SPLITS></RESULT><RESULT eventid="35" heatid="373" lane="2" points="308" resultid="2776" swimtime="00:00:36.14"><SPLITS/></RESULT><RESULT eventid="39" heatid="441" lane="6" points="400" resultid="3294" swimtime="00:01:10.13"><SPLITS><SPLIT distance="50" swimtime="00:00:32.97"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="349" birthdate="2010-01-01" firstname="Marie" gender="F" lastname="Starklauf" license="406868"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="48" lane="8" points="329" resultid="366" swimtime="00:05:42.39"><SPLITS><SPLIT distance="100" swimtime="00:01:15.64"/><SPLIT distance="200" swimtime="00:02:42.17"/><SPLIT distance="300" swimtime="00:04:13.03"/></SPLITS></RESULT><RESULT eventid="7" heatid="90" lane="3" points="410" resultid="675" swimtime="00:03:06.91"><SPLITS><SPLIT distance="50" swimtime="00:00:40.10"/><SPLIT distance="100" swimtime="00:01:27.70"/><SPLIT distance="150" swimtime="00:02:18.24"/></SPLITS></RESULT><RESULT eventid="17" heatid="230" lane="5" points="342" resultid="1736" swimtime="00:11:32.79"><SPLITS><SPLIT distance="100" swimtime="00:01:19.62"/><SPLIT distance="200" swimtime="00:02:46.71"/><SPLIT distance="300" swimtime="00:04:14.99"/><SPLIT distance="400" swimtime="00:05:43.83"/><SPLIT distance="500" swimtime="00:07:11.92"/><SPLIT distance="600" swimtime="00:08:39.83"/><SPLIT distance="700" swimtime="00:10:08.42"/></SPLITS></RESULT><RESULT eventid="31" heatid="343" lane="6" points="484" resultid="2560" swimtime="00:01:21.63"><SPLITS><SPLIT distance="50" swimtime="00:00:37.54"/></SPLITS></RESULT><RESULT eventid="37" heatid="407" lane="8" points="322" resultid="3038" swimtime="00:02:59.83"><SPLITS><SPLIT distance="50" swimtime="00:00:43.79"/><SPLIT distance="100" swimtime="00:01:28.94"/><SPLIT distance="150" swimtime="00:02:16.00"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="351" birthdate="2013-01-01" firstname="Marie" gender="F" lastname="Schellenberger" license="444718"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="49" lane="2" points="389" resultid="368" swimtime="00:05:23.84"><SPLITS><SPLIT distance="100" swimtime="00:01:15.06"/><SPLIT distance="200" swimtime="00:02:38.17"/><SPLIT distance="300" swimtime="00:04:01.84"/></SPLITS></RESULT><RESULT eventid="7" heatid="89" lane="4" points="406" resultid="668" swimtime="00:03:07.51"><SPLITS><SPLIT distance="50" swimtime="00:00:43.46"/><SPLIT distance="100" swimtime="00:01:32.24"/><SPLIT distance="150" swimtime="00:02:20.61"/></SPLITS></RESULT><RESULT eventid="11" heatid="169" lane="3" points="397" resultid="1277" swimtime="00:02:51.47"><SPLITS><SPLIT distance="50" swimtime="00:00:39.68"/><SPLIT distance="100" swimtime="00:01:25.19"/><SPLIT distance="150" swimtime="00:02:12.43"/></SPLITS></RESULT><RESULT eventid="25" heatid="248" lane="4" resultid="1840" swimtime="00:00:47.66"><SPLITS/></RESULT><RESULT eventid="31" heatid="341" lane="6" points="412" resultid="2544" swimtime="00:01:26.18"><SPLITS><SPLIT distance="50" swimtime="00:00:40.89"/></SPLITS></RESULT><RESULT eventid="35" heatid="373" lane="7" points="287" resultid="2781" swimtime="00:00:37.01"><SPLITS/></RESULT><RESULT eventid="39" heatid="440" lane="1" points="395" resultid="3282" swimtime="00:01:10.45"><SPLITS><SPLIT distance="50" swimtime="00:00:34.23"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="390" birthdate="2013-01-01" firstname="Joshua" gender="M" lastname="Baumüller" license="457275"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="55" lane="4" points="195" resultid="413" swimtime="00:06:19.28"><SPLITS><SPLIT distance="100" swimtime="00:01:24.96"/><SPLIT distance="200" swimtime="00:03:03.07"/><SPLIT distance="300" swimtime="00:04:43.89"/></SPLITS></RESULT><RESULT eventid="8" heatid="95" lane="8" points="151" resultid="717" swimtime="00:03:56.31"><SPLITS><SPLIT distance="50" swimtime="00:00:51.96"/><SPLIT distance="100" swimtime="00:01:51.67"/><SPLIT distance="150" swimtime="00:02:55.50"/></SPLITS></RESULT><RESULT eventid="10" heatid="138" lane="4" points="183" resultid="1040" swimtime="00:00:36.77"><SPLITS/></RESULT><RESULT eventid="12" heatid="177" lane="7" points="149" resultid="1341" swimtime="00:03:34.63"><SPLITS><SPLIT distance="50" swimtime="00:00:50.55"/><SPLIT distance="100" swimtime="00:01:46.26"/><SPLIT distance="150" swimtime="00:02:46.62"/></SPLITS></RESULT><RESULT eventid="24" heatid="245" lane="2" resultid="1821" swimtime="00:01:00.53"><SPLITS/></RESULT><RESULT eventid="30" heatid="313" lane="5" points="179" resultid="2331" swimtime="00:03:00.96"><SPLITS><SPLIT distance="50" swimtime="00:00:40.24"/><SPLIT distance="100" swimtime="00:01:27.06"/><SPLIT distance="150" swimtime="00:02:16.33"/></SPLITS></RESULT><RESULT eventid="36" heatid="386" lane="2" points="115" resultid="2872" swimtime="00:00:45.75"><SPLITS/></RESULT><RESULT eventid="40" heatid="459" lane="6" points="189" resultid="3434" swimtime="00:01:21.65"><SPLITS><SPLIT distance="50" swimtime="00:00:39.04"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="391" birthdate="2013-01-01" firstname="Aeneas" gender="M" lastname="Lange" license="450217"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="55" lane="5" points="161" resultid="414" swimtime="00:06:44.11"><SPLITS><SPLIT distance="100" swimtime="00:01:28.36"/><SPLIT distance="200" swimtime="00:03:11.28"/><SPLIT distance="300" swimtime="00:04:57.28"/></SPLITS></RESULT><RESULT eventid="6" heatid="72" lane="4" points="81" resultid="539" swimtime="00:01:53.90"><SPLITS><SPLIT distance="50" swimtime="00:00:49.76"/></SPLITS></RESULT><RESULT eventid="10" heatid="141" lane="5" points="161" resultid="1063" swimtime="00:00:38.40"><SPLITS/></RESULT><RESULT eventid="12" heatid="176" lane="7" points="126" resultid="1334" swimtime="00:03:47.31"><SPLITS><SPLIT distance="50" swimtime="00:00:50.45"/><SPLIT distance="100" swimtime="00:01:50.63"/><SPLIT distance="150" swimtime="00:02:55.64"/></SPLITS></RESULT><RESULT eventid="24" heatid="245" lane="1" resultid="1820" swimtime="00:00:58.39"><SPLITS/></RESULT><RESULT eventid="30" heatid="310" lane="4" points="153" resultid="2307" swimtime="00:03:10.46"><SPLITS><SPLIT distance="50" swimtime="00:00:38.52"/><SPLIT distance="100" swimtime="00:01:27.51"/><SPLIT distance="150" swimtime="00:02:18.40"/></SPLITS></RESULT><RESULT eventid="36" heatid="386" lane="5" points="105" resultid="2875" swimtime="00:00:47.11"><SPLITS/></RESULT><RESULT eventid="40" heatid="458" lane="2" points="165" resultid="3422" swimtime="00:01:25.40"><SPLITS><SPLIT distance="50" swimtime="00:00:38.96"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="403" birthdate="2010-01-01" firstname="Leo" gender="M" lastname="Gebhard" license="425301"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="57" lane="4" points="302" resultid="429" swimtime="00:05:27.78"><SPLITS><SPLIT distance="100" swimtime="00:01:12.57"/><SPLIT distance="200" swimtime="00:02:37.82"/><SPLIT distance="300" swimtime="00:04:04.78"/></SPLITS></RESULT><RESULT eventid="6" heatid="75" lane="7" points="197" resultid="565" swimtime="00:01:24.94"><SPLITS><SPLIT distance="50" swimtime="00:00:37.80"/></SPLITS></RESULT><RESULT eventid="10" heatid="148" lane="7" points="355" resultid="1120" swimtime="00:00:29.51"><SPLITS/></RESULT><RESULT eventid="12" heatid="183" lane="3" points="293" resultid="1384" swimtime="00:02:51.46"><SPLITS><SPLIT distance="50" swimtime="00:00:38.95"/><SPLIT distance="100" swimtime="00:01:23.41"/><SPLIT distance="150" swimtime="00:02:14.09"/></SPLITS></RESULT><RESULT eventid="30" heatid="317" lane="7" points="324" resultid="2364" swimtime="00:02:28.39"><SPLITS><SPLIT distance="50" swimtime="00:00:32.57"/><SPLIT distance="100" swimtime="00:01:09.50"/><SPLIT distance="150" swimtime="00:01:48.98"/></SPLITS></RESULT><RESULT eventid="36" heatid="392" lane="1" points="256" resultid="2918" swimtime="00:00:35.05"><SPLITS/></RESULT><RESULT eventid="40" heatid="467" lane="2" points="354" resultid="3492" swimtime="00:01:06.19"><SPLITS><SPLIT distance="50" swimtime="00:00:31.41"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="405" birthdate="2012-01-01" firstname="Nils" gender="M" lastname="Wöhner" license="437511"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="57" lane="7" points="284" resultid="432" swimtime="00:05:34.58"><SPLITS><SPLIT distance="100" swimtime="00:01:18.53"/><SPLIT distance="200" swimtime="00:02:45.12"/><SPLIT distance="300" swimtime="00:04:12.13"/></SPLITS></RESULT><RESULT eventid="6" heatid="74" lane="4" points="171" resultid="554" swimtime="00:01:29.06"><SPLITS><SPLIT distance="50" swimtime="00:00:39.40"/></SPLITS></RESULT><RESULT eventid="10" heatid="145" lane="6" points="258" resultid="1095" swimtime="00:00:32.82"><SPLITS/></RESULT><RESULT eventid="12" heatid="181" lane="6" points="226" resultid="1371" swimtime="00:03:06.89"><SPLITS><SPLIT distance="50" swimtime="00:00:41.87"/><SPLIT distance="100" swimtime="00:01:31.20"/><SPLIT distance="150" swimtime="00:02:28.94"/></SPLITS></RESULT><RESULT eventid="28" heatid="283" lane="1" points="216" resultid="2101" swimtime="00:00:39.46"><SPLITS/></RESULT><RESULT eventid="30" heatid="319" lane="4" points="284" resultid="2377" swimtime="00:02:35.00"><SPLITS><SPLIT distance="50" swimtime="00:00:35.67"/><SPLIT distance="100" swimtime="00:01:15.89"/><SPLIT distance="150" swimtime="00:01:56.25"/></SPLITS></RESULT><RESULT eventid="36" heatid="391" lane="2" points="197" resultid="2911" swimtime="00:00:38.23"><SPLITS/></RESULT><RESULT eventid="40" heatid="465" lane="2" points="275" resultid="3476" swimtime="00:01:12.05"><SPLITS><SPLIT distance="50" swimtime="00:00:34.53"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="409" birthdate="2013-01-01" firstname="Hendrik" gender="M" lastname="Schick" license="447027"><HANDICAP/><ENTRIES/><RESULTS><RESULT comment="10:58 Start vor dem Startsignal" eventid="4" heatid="58" lane="5" resultid="438" status="DSQ" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="12" heatid="182" lane="4" points="282" resultid="1377" swimtime="00:02:53.70"><SPLITS><SPLIT distance="50" swimtime="00:00:37.32"/><SPLIT distance="100" swimtime="00:01:22.62"/><SPLIT distance="150" swimtime="00:02:16.14"/></SPLITS></RESULT><RESULT eventid="14" heatid="221" lane="2" points="260" resultid="1675" swimtime="00:01:20.78"><SPLITS><SPLIT distance="50" swimtime="00:00:39.45"/></SPLITS></RESULT><RESULT eventid="24" heatid="245" lane="4" resultid="1823" swimtime="00:00:47.05"><SPLITS/></RESULT><RESULT eventid="28" heatid="281" lane="5" points="232" resultid="2089" swimtime="00:00:38.58"><SPLITS/></RESULT><RESULT eventid="30" heatid="319" lane="5" points="293" resultid="2378" swimtime="00:02:33.48"><SPLITS><SPLIT distance="50" swimtime="00:00:35.55"/><SPLIT distance="100" swimtime="00:01:15.50"/><SPLIT distance="150" swimtime="00:01:55.44"/></SPLITS></RESULT><RESULT eventid="38" heatid="417" lane="3" points="285" resultid="3109" swimtime="00:02:49.91"><SPLITS><SPLIT distance="50" swimtime="00:00:40.57"/><SPLIT distance="100" swimtime="00:01:24.02"/><SPLIT distance="150" swimtime="00:02:09.00"/></SPLITS></RESULT><RESULT eventid="40" heatid="465" lane="5" points="283" resultid="3479" swimtime="00:01:11.36"><SPLITS><SPLIT distance="50" swimtime="00:00:34.53"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="438" birthdate="2009-01-01" firstname="Samuel" gender="M" lastname="Lang" license="392828"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="62" lane="8" points="556" resultid="468" swimtime="00:04:27.63"><SPLITS><SPLIT distance="100" swimtime="00:01:02.79"/><SPLIT distance="200" swimtime="00:02:09.87"/><SPLIT distance="300" swimtime="00:03:18.19"/></SPLITS></RESULT><RESULT eventid="6" heatid="79" lane="8" points="466" resultid="597" swimtime="00:01:03.74"><SPLITS><SPLIT distance="50" swimtime="00:00:30.24"/></SPLITS></RESULT><RESULT eventid="10" heatid="153" lane="1" points="478" resultid="1154" swimtime="00:00:26.74"><SPLITS/></RESULT><RESULT eventid="30" heatid="325" lane="1" points="575" resultid="2419" swimtime="00:02:02.60"><SPLITS><SPLIT distance="50" swimtime="00:00:28.59"/><SPLIT distance="100" swimtime="00:00:59.41"/><SPLIT distance="150" swimtime="00:01:30.96"/></SPLITS></RESULT><RESULT eventid="34" heatid="362" lane="5" points="502" resultid="2693" swimtime="00:02:18.76"><SPLITS><SPLIT distance="50" swimtime="00:00:29.54"/><SPLIT distance="100" swimtime="00:01:05.24"/><SPLIT distance="150" swimtime="00:01:42.50"/></SPLITS></RESULT><RESULT eventid="36" heatid="398" lane="8" points="468" resultid="2973" swimtime="00:00:28.67"><SPLITS/></RESULT><RESULT eventid="40" heatid="472" lane="2" points="576" resultid="3531" swimtime="00:00:56.29"><SPLITS><SPLIT distance="50" swimtime="00:00:26.74"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="446" birthdate="2011-01-01" firstname="Charlotte" gender="F" lastname="Hammann" license="423699"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="5" heatid="65" lane="5" points="265" resultid="485" swimtime="00:01:26.32"><SPLITS><SPLIT distance="50" swimtime="00:00:38.89"/></SPLITS></RESULT><RESULT eventid="11" heatid="166" lane="7" points="334" resultid="1257" swimtime="00:03:01.71"><SPLITS><SPLIT distance="50" swimtime="00:00:39.62"/><SPLIT distance="100" swimtime="00:01:24.36"/><SPLIT distance="150" swimtime="00:02:17.63"/></SPLITS></RESULT><RESULT eventid="13" heatid="206" lane="5" points="346" resultid="1564" swimtime="00:01:21.78"><SPLITS><SPLIT distance="50" swimtime="00:00:40.86"/></SPLITS></RESULT><RESULT eventid="27" heatid="269" lane="7" points="416" resultid="2001" swimtime="00:00:36.14"><SPLITS/></RESULT><RESULT eventid="35" heatid="376" lane="2" points="304" resultid="2799" swimtime="00:00:36.33"><SPLITS/></RESULT><RESULT eventid="37" heatid="409" lane="8" points="328" resultid="3054" swimtime="00:02:58.86"><SPLITS><SPLIT distance="50" swimtime="00:00:42.60"/><SPLIT distance="100" swimtime="00:01:27.19"/><SPLIT distance="150" swimtime="00:02:14.97"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="449" birthdate="2011-01-01" firstname="Olivia" gender="F" lastname="Lang" license="425304"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="5" heatid="66" lane="6" points="295" resultid="494" swimtime="00:01:23.25"><SPLITS><SPLIT distance="50" swimtime="00:00:37.50"/></SPLITS></RESULT><RESULT eventid="9" heatid="123" lane="8" points="364" resultid="935" swimtime="00:00:33.14"><SPLITS/></RESULT><RESULT eventid="11" heatid="165" lane="5" points="328" resultid="1247" swimtime="00:03:02.81"><SPLITS><SPLIT distance="50" swimtime="00:00:40.25"/><SPLIT distance="100" swimtime="00:01:29.02"/><SPLIT distance="150" swimtime="00:02:23.48"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="492" birthdate="2010-01-01" firstname="Jannik" gender="M" lastname="Hünniger" license="409224"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="6" heatid="78" lane="2" points="425" resultid="583" swimtime="00:01:05.77"><SPLITS><SPLIT distance="50" swimtime="00:00:30.33"/></SPLITS></RESULT><RESULT eventid="10" heatid="155" lane="4" points="553" resultid="1172" swimtime="00:00:25.47"><SPLITS/></RESULT><RESULT eventid="14" heatid="224" lane="6" points="429" resultid="1702" swimtime="00:01:08.39"><SPLITS><SPLIT distance="50" swimtime="00:00:31.97"/></SPLITS></RESULT><RESULT eventid="30" heatid="323" lane="5" points="462" resultid="2407" swimtime="00:02:11.93"><SPLITS><SPLIT distance="50" swimtime="00:00:29.20"/><SPLIT distance="100" swimtime="00:01:03.08"/><SPLIT distance="150" swimtime="00:01:38.46"/></SPLITS></RESULT><RESULT eventid="40" heatid="472" lane="4" points="513" resultid="3533" swimtime="00:00:58.50"><SPLITS><SPLIT distance="50" swimtime="00:00:28.07"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="509" birthdate="2009-01-01" firstname="Greta" gender="F" lastname="Lange" license="377374"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="7" heatid="91" lane="5" points="477" resultid="685" swimtime="00:02:57.82"><SPLITS><SPLIT distance="50" swimtime="00:00:40.20"/><SPLIT distance="100" swimtime="00:01:25.61"/><SPLIT distance="150" swimtime="00:02:11.49"/></SPLITS></RESULT><RESULT eventid="9" heatid="127" lane="3" points="412" resultid="961" swimtime="00:00:31.79"><SPLITS/></RESULT><RESULT eventid="31" heatid="342" lane="3" points="444" resultid="2549" swimtime="00:01:24.03"><SPLITS><SPLIT distance="50" swimtime="00:00:40.06"/></SPLITS></RESULT><RESULT eventid="35" heatid="376" lane="8" points="320" resultid="2805" swimtime="00:00:35.68"><SPLITS/></RESULT><RESULT eventid="39" heatid="444" lane="4" points="413" resultid="3316" swimtime="00:01:09.41"><SPLITS><SPLIT distance="50" swimtime="00:00:32.73"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="515" birthdate="2016-01-01" firstname="Lotte" gender="F" lastname="Fankel" license="454670"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="9" heatid="110" lane="2" points="275" resultid="826" swimtime="00:00:36.38"><SPLITS/></RESULT><RESULT eventid="13" heatid="196" lane="7" points="204" resultid="1486" swimtime="00:01:37.57"><SPLITS><SPLIT distance="50" swimtime="00:00:47.42"/></SPLITS></RESULT><RESULT eventid="27" heatid="258" lane="3" points="180" resultid="1910" swimtime="00:00:47.77"><SPLITS/></RESULT><RESULT eventid="29" heatid="293" lane="5" points="247" resultid="2178" swimtime="00:02:59.85"><SPLITS><SPLIT distance="50" swimtime="00:00:41.88"/><SPLIT distance="100" swimtime="00:01:28.11"/><SPLIT distance="150" swimtime="00:02:15.79"/></SPLITS></RESULT><RESULT eventid="35" heatid="366" lane="7" points="129" resultid="2725" swimtime="00:00:48.28"><SPLITS/></RESULT><RESULT eventid="37" heatid="403" lane="7" points="222" resultid="3005" swimtime="00:03:23.62"><SPLITS><SPLIT distance="50" swimtime="00:00:48.72"/><SPLIT distance="100" swimtime="00:01:40.72"/><SPLIT distance="150" swimtime="00:02:34.31"/></SPLITS></RESULT><RESULT eventid="39" heatid="430" lane="2" points="256" resultid="3203" swimtime="00:01:21.41"><SPLITS><SPLIT distance="50" swimtime="00:00:39.39"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="533" birthdate="2010-01-01" firstname="Clara" gender="F" lastname="Ehrlich" license="406861"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="9" heatid="130" lane="4" points="544" resultid="986" swimtime="00:00:28.98"><SPLITS/></RESULT><RESULT eventid="13" heatid="208" lane="2" points="515" resultid="1576" swimtime="00:01:11.65"><SPLITS><SPLIT distance="50" swimtime="00:00:34.32"/></SPLITS></RESULT><RESULT eventid="27" heatid="272" lane="1" points="478" resultid="2018" swimtime="00:00:34.50"><SPLITS/></RESULT><RESULT eventid="37" heatid="412" lane="1" points="492" resultid="3071" swimtime="00:02:36.23"><SPLITS><SPLIT distance="100" swimtime="00:01:13.94"/></SPLITS></RESULT><RESULT eventid="39" heatid="449" lane="2" points="517" resultid="3352" swimtime="00:01:04.39"><SPLITS><SPLIT distance="50" swimtime="00:00:30.46"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="548" birthdate="2014-01-01" firstname="Mika" gender="M" lastname="Fankel" license="454669"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="10" heatid="145" lane="3" points="249" resultid="1092" swimtime="00:00:33.23"><SPLITS/></RESULT><RESULT eventid="12" heatid="183" lane="2" points="272" resultid="1383" swimtime="00:02:55.82"><SPLITS><SPLIT distance="50" swimtime="00:00:37.76"/><SPLIT distance="100" swimtime="00:01:23.02"/><SPLIT distance="150" swimtime="00:02:16.75"/></SPLITS></RESULT><RESULT eventid="14" heatid="220" lane="6" points="227" resultid="1671" swimtime="00:01:24.55"><SPLITS><SPLIT distance="50" swimtime="00:00:40.81"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="556" birthdate="2011-01-01" firstname="Bartosz" gender="M" lastname="Gorczynski" license="429037"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="10" heatid="153" lane="7" points="483" resultid="1160" swimtime="00:00:26.64"><SPLITS/></RESULT><RESULT eventid="12" heatid="188" lane="8" points="429" resultid="1427" swimtime="00:02:31.14"><SPLITS><SPLIT distance="50" swimtime="00:00:31.76"/><SPLIT distance="100" swimtime="00:01:12.37"/><SPLIT distance="150" swimtime="00:01:57.58"/></SPLITS></RESULT><RESULT eventid="28" heatid="284" lane="2" points="420" resultid="2110" swimtime="00:00:31.66"><SPLITS/></RESULT><RESULT eventid="36" heatid="396" lane="8" points="411" resultid="2957" swimtime="00:00:29.94"><SPLITS/></RESULT><RESULT eventid="40" heatid="472" lane="8" points="495" resultid="3537" swimtime="00:00:59.22"><SPLITS><SPLIT distance="50" swimtime="00:00:28.47"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="602" birthdate="2012-01-01" firstname="Ferdinand" gender="M" lastname="Behrens" license="457278"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="30" heatid="312" lane="3" points="209" resultid="2321" swimtime="00:02:51.86"><SPLITS><SPLIT distance="50" swimtime="00:00:36.04"/><SPLIT distance="100" swimtime="00:01:20.29"/><SPLIT distance="150" swimtime="00:02:08.22"/></SPLITS></RESULT><RESULT eventid="32" heatid="350" lane="4" points="201" resultid="2608" swimtime="00:01:37.06"><SPLITS><SPLIT distance="50" swimtime="00:00:43.54"/></SPLITS></RESULT><RESULT eventid="36" heatid="385" lane="6" points="158" resultid="2868" swimtime="00:00:41.12"><SPLITS/></RESULT><RESULT eventid="40" heatid="459" lane="7" points="226" resultid="3435" swimtime="00:01:16.83"><SPLITS><SPLIT distance="50" swimtime="00:00:35.96"/></SPLITS></RESULT></RESULTS></ATHLETE></ATHLETES><RELAYS/></CLUB><CLUB name="Kinder- und Jugendschule &quot;Schkid&quot;" nation="UKR" shortname="Schkid" type="CLUB"><CONTACT city="Browary" country="UKR" name="Karolina Rusavska"/><OFFICIALS/><ATHLETES><ATHLETE athleteid="99" birthdate="2009-01-01" firstname="Sofiia" gender="F" lastname="Dotsenko"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="13" lane="7" points="161" resultid="99" swimtime="00:00:53.81"><SPLITS/></RESULT><RESULT eventid="9" heatid="113" lane="6" points="171" resultid="854" swimtime="00:00:42.61"><SPLITS/></RESULT><RESULT eventid="31" heatid="333" lane="1" points="162" resultid="2475" swimtime="00:01:57.54"><SPLITS><SPLIT distance="50" swimtime="00:00:55.68"/></SPLITS></RESULT><RESULT eventid="39" heatid="427" lane="1" points="158" resultid="3178" swimtime="00:01:35.65"><SPLITS><SPLIT distance="50" swimtime="00:00:43.65"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="270" birthdate="2011-01-01" firstname="Dmytro" gender="M" lastname="Dorogoi"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="36" lane="4" points="273" resultid="270" swimtime="00:00:39.98"><SPLITS/></RESULT><RESULT eventid="8" heatid="98" lane="3" points="272" resultid="736" swimtime="00:03:14.22"><SPLITS><SPLIT distance="50" swimtime="00:00:45.10"/><SPLIT distance="100" swimtime="00:01:36.29"/><SPLIT distance="150" swimtime="00:02:28.06"/></SPLITS></RESULT><RESULT eventid="12" heatid="179" lane="2" points="224" resultid="1351" swimtime="00:03:07.46"><SPLITS><SPLIT distance="50" swimtime="00:00:45.67"/><SPLIT distance="100" swimtime="00:01:36.73"/><SPLIT distance="150" swimtime="00:02:26.50"/></SPLITS></RESULT><RESULT eventid="32" heatid="352" lane="3" points="271" resultid="2622" swimtime="00:01:27.88"><SPLITS><SPLIT distance="50" swimtime="00:00:42.97"/></SPLITS></RESULT><RESULT eventid="40" heatid="463" lane="5" points="213" resultid="3463" swimtime="00:01:18.44"><SPLITS><SPLIT distance="50" swimtime="00:00:37.42"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="299" birthdate="2008-01-01" firstname="Myron" gender="M" lastname="Pinchuk"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="40" lane="1" points="534" resultid="299" swimtime="00:00:31.98"><SPLITS/></RESULT><RESULT eventid="8" heatid="101" lane="1" points="476" resultid="757" swimtime="00:02:41.29"><SPLITS><SPLIT distance="50" swimtime="00:00:37.95"/><SPLIT distance="100" swimtime="00:01:20.89"/><SPLIT distance="150" swimtime="00:02:01.80"/></SPLITS></RESULT><RESULT eventid="10" heatid="151" lane="1" points="447" resultid="1138" swimtime="00:00:27.33"><SPLITS/></RESULT><RESULT eventid="32" heatid="356" lane="7" points="498" resultid="2656" swimtime="00:01:11.73"><SPLITS><SPLIT distance="50" swimtime="00:00:32.87"/></SPLITS></RESULT><RESULT eventid="36" heatid="395" lane="4" points="416" resultid="2945" swimtime="00:00:29.82"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="333" birthdate="2010-01-01" firstname="Yelyzaveta" gender="F" lastname="Horban"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="45" lane="6" points="295" resultid="341" swimtime="00:05:55.10"><SPLITS><SPLIT distance="100" swimtime="00:01:21.92"/><SPLIT distance="200" swimtime="00:02:53.27"/><SPLIT distance="300" swimtime="00:04:26.95"/></SPLITS></RESULT><RESULT eventid="9" heatid="119" lane="1" points="320" resultid="896" swimtime="00:00:34.57"><SPLITS/></RESULT><RESULT eventid="29" heatid="299" lane="7" points="327" resultid="2228" swimtime="00:02:43.94"><SPLITS><SPLIT distance="50" swimtime="00:00:37.80"/><SPLIT distance="100" swimtime="00:01:20.24"/><SPLIT distance="150" swimtime="00:02:02.47"/></SPLITS></RESULT><RESULT eventid="39" heatid="439" lane="8" points="334" resultid="3281" swimtime="00:01:14.48"><SPLITS><SPLIT distance="50" swimtime="00:00:36.26"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="415" birthdate="2009-01-01" firstname="Oleksandr" gender="M" lastname="Mizin"><HANDICAP/><ENTRIES/><RESULTS><RESULT comment="11:07 Der Schwimmer hat bei Doppelbahnbelegung seine Bahnseite verlassen und den anderen Schwimmer behindert" eventid="4" heatid="59" lane="4" resultid="444" status="DSQ" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="12" heatid="186" lane="6" points="356" resultid="1409" swimtime="00:02:40.82"><SPLITS><SPLIT distance="50" swimtime="00:00:36.17"/><SPLIT distance="100" swimtime="00:01:19.03"/><SPLIT distance="150" swimtime="00:02:05.65"/></SPLITS></RESULT><RESULT eventid="30" heatid="321" lane="1" points="335" resultid="2390" swimtime="00:02:26.83"><SPLITS><SPLIT distance="50" swimtime="00:00:36.38"/><SPLIT distance="100" swimtime="00:01:14.58"/><SPLIT distance="150" swimtime="00:01:52.24"/></SPLITS></RESULT><RESULT eventid="42" heatid="479" lane="7" points="372" resultid="3583" swimtime="00:05:38.96"><SPLITS><SPLIT distance="50" swimtime="00:00:36.32"/><SPLIT distance="100" swimtime="00:01:20.68"/><SPLIT distance="150" swimtime="00:02:03.82"/><SPLIT distance="200" swimtime="00:02:45.92"/><SPLIT distance="250" swimtime="00:03:34.89"/><SPLIT distance="300" swimtime="00:04:24.66"/><SPLIT distance="350" swimtime="00:05:02.47"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="419" birthdate="2011-01-01" firstname="Vladyslav" gender="M" lastname="Usatiuk"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="59" lane="8" points="290" resultid="448" swimtime="00:05:32.41"><SPLITS><SPLIT distance="100" swimtime="00:01:16.63"/><SPLIT distance="200" swimtime="00:02:42.91"/><SPLIT distance="300" swimtime="00:04:09.20"/></SPLITS></RESULT><RESULT eventid="10" heatid="148" lane="2" points="274" resultid="1115" swimtime="00:00:32.17"><SPLITS/></RESULT><RESULT eventid="30" heatid="320" lane="1" points="291" resultid="2382" swimtime="00:02:33.80"><SPLITS><SPLIT distance="50" swimtime="00:00:35.69"/><SPLIT distance="100" swimtime="00:01:15.19"/><SPLIT distance="150" swimtime="00:01:55.67"/></SPLITS></RESULT><RESULT eventid="40" heatid="467" lane="5" points="321" resultid="3494" swimtime="00:01:08.37"><SPLITS><SPLIT distance="50" swimtime="00:00:32.96"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="443" birthdate="2012-01-01" firstname="Mariia" gender="F" lastname="Dotsenko"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="5" heatid="64" lane="8" points="156" resultid="480" swimtime="00:01:42.88"><SPLITS><SPLIT distance="50" swimtime="00:00:47.47"/></SPLITS></RESULT><RESULT comment="13:06 Die Sportlerin führte die Arme während der Schwimmstrecke nicht gleichzeitig über Wasser nach vorne" eventid="33" heatid="357" lane="5" resultid="2660" status="DSQ" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="35" heatid="367" lane="6" points="171" resultid="2732" swimtime="00:00:44.00"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="479" birthdate="2009-01-01" firstname="Anton" gender="M" lastname="Cherednychok"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="6" heatid="75" lane="2" points="227" resultid="560" swimtime="00:01:21.01"><SPLITS><SPLIT distance="50" swimtime="00:00:34.33"/></SPLITS></RESULT><RESULT eventid="10" heatid="153" lane="8" points="415" resultid="1161" swimtime="00:00:28.03"><SPLITS/></RESULT><RESULT eventid="30" heatid="318" lane="4" points="193" resultid="2369" swimtime="00:02:56.28"><SPLITS><SPLIT distance="50" swimtime="00:00:31.82"/><SPLIT distance="100" swimtime="00:01:11.21"/><SPLIT distance="150" swimtime="00:02:01.23"/></SPLITS></RESULT><RESULT eventid="36" heatid="394" lane="2" points="307" resultid="2935" swimtime="00:00:32.98"><SPLITS/></RESULT><RESULT eventid="40" heatid="470" lane="4" points="376" resultid="3517" swimtime="00:01:04.92"><SPLITS><SPLIT distance="50" swimtime="00:00:30.52"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="484" birthdate="2009-01-01" firstname="Yaroslav" gender="M" lastname="Chernikov"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="6" heatid="76" lane="3" points="383" resultid="569" swimtime="00:01:08.07"><SPLITS><SPLIT distance="50" swimtime="00:00:30.61"/></SPLITS></RESULT><RESULT eventid="14" heatid="223" lane="3" points="359" resultid="1692" swimtime="00:01:12.54"><SPLITS><SPLIT distance="50" swimtime="00:00:36.03"/></SPLITS></RESULT><RESULT eventid="28" heatid="285" lane="2" resultid="2117" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="36" heatid="397" lane="1" points="431" resultid="2958" swimtime="00:00:29.47"><SPLITS/></RESULT><RESULT eventid="42" heatid="479" lane="6" points="369" resultid="3582" swimtime="00:05:39.86"><SPLITS><SPLIT distance="50" swimtime="00:00:32.17"/><SPLIT distance="100" swimtime="00:01:11.16"/><SPLIT distance="150" swimtime="00:01:54.97"/><SPLIT distance="200" swimtime="00:02:36.61"/><SPLIT distance="250" swimtime="00:03:27.26"/><SPLIT distance="300" swimtime="00:04:18.48"/><SPLIT distance="350" swimtime="00:05:01.47"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="494" birthdate="2009-01-01" firstname="Yehor" gender="M" lastname="Ishenko"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="6" heatid="78" lane="4" points="511" resultid="585" swimtime="00:01:01.82"><SPLITS><SPLIT distance="50" swimtime="00:00:27.51"/></SPLITS></RESULT><RESULT eventid="10" heatid="157" lane="8" points="528" resultid="1191" swimtime="00:00:25.86"><SPLITS/></RESULT><RESULT eventid="14" heatid="224" lane="5" points="498" resultid="1701" swimtime="00:01:05.09"><SPLITS><SPLIT distance="50" swimtime="00:00:31.15"/></SPLITS></RESULT><RESULT eventid="28" heatid="287" lane="1" points="462" resultid="2132" swimtime="00:00:30.66"><SPLITS/></RESULT><RESULT eventid="36" heatid="400" lane="8" points="532" resultid="2988" swimtime="00:00:27.48"><SPLITS/></RESULT><RESULT eventid="40" heatid="474" lane="4" points="576" resultid="3548" swimtime="00:00:56.30"><SPLITS><SPLIT distance="50" swimtime="00:00:27.25"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="524" birthdate="2009-01-01" firstname="Dariia" gender="F" lastname="Tsyts"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="9" heatid="123" lane="4" points="424" resultid="931" swimtime="00:00:31.49"><SPLITS/></RESULT><RESULT eventid="11" heatid="166" lane="4" points="325" resultid="1254" swimtime="00:03:03.28"><SPLITS><SPLIT distance="50" swimtime="00:00:38.08"/><SPLIT distance="100" swimtime="00:01:27.54"/><SPLIT distance="150" swimtime="00:02:21.06"/></SPLITS></RESULT><RESULT eventid="29" heatid="294" lane="2" points="309" resultid="2183" swimtime="00:02:46.94"><SPLITS><SPLIT distance="50" swimtime="00:00:36.23"/><SPLIT distance="100" swimtime="00:01:17.82"/><SPLIT distance="150" swimtime="00:02:03.22"/></SPLITS></RESULT><RESULT eventid="39" heatid="442" lane="1" points="380" resultid="3297" swimtime="00:01:11.37"><SPLITS><SPLIT distance="50" swimtime="00:00:33.64"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="546" birthdate="2011-01-01" firstname="Ihor" gender="M" lastname="Petrov"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="10" heatid="142" lane="2" points="182" resultid="1068" swimtime="00:00:36.85"><SPLITS/></RESULT><RESULT eventid="14" heatid="217" lane="5" points="161" resultid="1647" swimtime="00:01:34.66"><SPLITS><SPLIT distance="50" swimtime="00:00:45.12"/></SPLITS></RESULT><RESULT eventid="28" heatid="282" lane="8" points="163" resultid="2100" swimtime="00:00:43.36"><SPLITS/></RESULT><RESULT eventid="30" heatid="313" lane="4" points="152" resultid="2330" swimtime="00:03:10.88"><SPLITS><SPLIT distance="50" swimtime="00:00:41.70"/><SPLIT distance="100" swimtime="00:01:32.47"/><SPLIT distance="150" swimtime="00:02:22.52"/></SPLITS></RESULT><RESULT eventid="40" heatid="459" lane="3" points="166" resultid="3431" swimtime="00:01:25.15"><SPLITS><SPLIT distance="50" swimtime="00:00:41.10"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="563" birthdate="2010-01-01" firstname="Artem" gender="M" lastname="Musatenko"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="12" heatid="181" lane="1" points="229" resultid="1366" swimtime="00:03:06.24"><SPLITS><SPLIT distance="50" swimtime="00:00:37.75"/><SPLIT distance="100" swimtime="00:01:21.90"/><SPLIT distance="150" swimtime="00:02:18.82"/></SPLITS></RESULT><RESULT eventid="14" heatid="221" lane="7" points="254" resultid="1680" swimtime="00:01:21.43"><SPLITS><SPLIT distance="50" swimtime="00:00:39.20"/></SPLITS></RESULT><RESULT eventid="28" heatid="283" lane="2" points="263" resultid="2102" swimtime="00:00:36.97"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="564" birthdate="2011-01-01" firstname="Ivan" gender="M" lastname="Rusin"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="12" heatid="187" lane="5" points="223" resultid="1416" swimtime="00:03:07.94"><SPLITS><SPLIT distance="50" swimtime="00:00:39.32"/><SPLIT distance="100" swimtime="00:01:27.34"/><SPLIT distance="150" swimtime="00:02:26.30"/></SPLITS></RESULT><RESULT eventid="30" heatid="318" lane="5" points="238" resultid="2370" swimtime="00:02:44.55"><SPLITS><SPLIT distance="50" swimtime="00:00:36.25"/><SPLIT distance="100" swimtime="00:01:18.78"/><SPLIT distance="150" swimtime="00:02:01.81"/></SPLITS></RESULT><RESULT eventid="36" heatid="393" lane="8" points="206" resultid="2933" swimtime="00:00:37.65"><SPLITS/></RESULT><RESULT eventid="40" heatid="466" lane="3" points="275" resultid="3485" swimtime="00:01:11.99"><SPLITS><SPLIT distance="50" swimtime="00:00:34.44"/></SPLITS></RESULT></RESULTS></ATHLETE></ATHLETES><RELAYS><RELAY agemax="-1" agemin="-1" agetotalmax="14" agetotalmin="14" gender="M" name="1. Mannschaft" number="1"><ENTRIES/><RESULTS><RESULT eventid="44" heatid="483" lane="6" points="356" resultid="3599" swimtime="00:09:50.11"><SPLITS><SPLIT distance="50" swimtime="00:00:36.07"/><SPLIT distance="100" swimtime="00:01:15.56"/><SPLIT distance="150" swimtime="00:01:53.99"/><SPLIT distance="200" swimtime="00:02:30.39"/><SPLIT distance="250" swimtime="00:03:05.16"/><SPLIT distance="300" swimtime="00:03:46.18"/><SPLIT distance="350" swimtime="00:04:28.18"/><SPLIT distance="400" swimtime="00:05:07.48"/><SPLIT distance="450" swimtime="00:05:41.90"/><SPLIT distance="500" swimtime="00:06:21.60"/><SPLIT distance="550" swimtime="00:07:00.90"/><SPLIT distance="600" swimtime="00:07:39.80"/><SPLIT distance="650" swimtime="00:08:09.41"/><SPLIT distance="700" swimtime="00:08:42.79"/><SPLIT distance="750" swimtime="00:09:17.65"/></SPLITS><RELAYPOSITIONS><RELAYPOSITION athleteid="415" number="1"/><RELAYPOSITION athleteid="484" number="2"/><RELAYPOSITION athleteid="419" number="3"/><RELAYPOSITION athleteid="494" number="4"/></RELAYPOSITIONS></RESULT></RESULTS></RELAY></RELAYS></CLUB><CLUB code="4357" name="SV Grafing-Ebersberg" nation="GER" region="02" shortname="Grafing" type="CLUB"><CONTACT city="Haar" email="wettkampf.svge@googlemail.com" name="Hable, Sabrina" phone="08093 / 9444" street="Am Seestall 23" zip="85625"/><OFFICIALS/><ATHLETES><ATHLETE athleteid="105" birthdate="2014-01-01" firstname="Sophia" gender="F" lastname="Dörrer" license="477865"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="14" lane="5" points="265" resultid="105" swimtime="00:00:45.56"><SPLITS/></RESULT><RESULT eventid="7" heatid="83" lane="7" points="232" resultid="624" swimtime="00:03:45.84"><SPLITS><SPLIT distance="50" swimtime="00:00:49.93"/><SPLIT distance="100" swimtime="00:01:48.01"/><SPLIT distance="150" swimtime="00:02:47.11"/></SPLITS></RESULT><RESULT eventid="9" heatid="115" lane="4" points="307" resultid="868" swimtime="00:00:35.08"><SPLITS/></RESULT><RESULT eventid="11" heatid="158" lane="3" points="217" resultid="1192" swimtime="00:03:29.70"><SPLITS><SPLIT distance="50" swimtime="00:00:44.40"/><SPLIT distance="100" swimtime="00:01:41.31"/><SPLIT distance="150" swimtime="00:02:42.00"/></SPLITS></RESULT><RESULT eventid="31" heatid="336" lane="8" points="252" resultid="2506" swimtime="00:01:41.48"><SPLITS><SPLIT distance="50" swimtime="00:00:47.99"/></SPLITS></RESULT><RESULT eventid="37" heatid="402" lane="2" points="228" resultid="2993" swimtime="00:03:21.89"><SPLITS><SPLIT distance="50" swimtime="00:00:47.57"/><SPLIT distance="100" swimtime="00:01:40.32"/><SPLIT distance="150" swimtime="00:02:33.22"/></SPLITS></RESULT><RESULT eventid="39" heatid="428" lane="1" points="245" resultid="3186" swimtime="00:01:22.58"><SPLITS><SPLIT distance="50" swimtime="00:00:39.33"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="110" birthdate="2013-01-01" firstname="Felicia" gender="F" lastname="Lampl" license="466176"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="15" lane="2" points="242" resultid="110" swimtime="00:00:46.97"><SPLITS/></RESULT><RESULT eventid="7" heatid="85" lane="4" points="261" resultid="636" swimtime="00:03:37.34"><SPLITS><SPLIT distance="50" swimtime="00:00:49.02"/><SPLIT distance="100" swimtime="00:01:47.02"/><SPLIT distance="150" swimtime="00:02:43.25"/></SPLITS></RESULT><RESULT eventid="9" heatid="114" lane="8" points="238" resultid="864" swimtime="00:00:38.17"><SPLITS/></RESULT><RESULT eventid="27" heatid="261" lane="3" points="231" resultid="1934" swimtime="00:00:43.96"><SPLITS/></RESULT><RESULT eventid="31" heatid="336" lane="7" points="277" resultid="2505" swimtime="00:01:38.29"><SPLITS><SPLIT distance="50" swimtime="00:00:46.43"/></SPLITS></RESULT><RESULT eventid="39" heatid="429" lane="2" points="218" resultid="3195" swimtime="00:01:25.81"><SPLITS><SPLIT distance="50" swimtime="00:00:40.57"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="137" birthdate="2007-01-01" firstname="Lisa" gender="F" lastname="Blankenburg" license="368541"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="18" lane="5" points="251" resultid="137" swimtime="00:00:46.39"><SPLITS/></RESULT><RESULT eventid="7" heatid="87" lane="5" points="287" resultid="653" swimtime="00:03:30.47"><SPLITS><SPLIT distance="50" swimtime="00:00:45.62"/><SPLIT distance="100" swimtime="00:01:38.09"/><SPLIT distance="150" swimtime="00:02:34.44"/></SPLITS></RESULT><RESULT eventid="9" heatid="116" lane="6" points="257" resultid="878" swimtime="00:00:37.20"><SPLITS/></RESULT><RESULT eventid="29" heatid="297" lane="2" points="278" resultid="2207" swimtime="00:02:52.93"><SPLITS><SPLIT distance="50" swimtime="00:00:38.53"/><SPLIT distance="100" swimtime="00:01:21.66"/><SPLIT distance="150" swimtime="00:02:08.77"/></SPLITS></RESULT><RESULT eventid="31" heatid="338" lane="2" points="295" resultid="2516" swimtime="00:01:36.24"><SPLITS><SPLIT distance="50" swimtime="00:00:45.91"/></SPLITS></RESULT><RESULT eventid="39" heatid="435" lane="6" points="237" resultid="3247" swimtime="00:01:23.48"><SPLITS><SPLIT distance="50" swimtime="00:00:38.72"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="142" birthdate="2009-01-01" firstname="Sarah" gender="F" lastname="Lechleiter" license="423199"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="19" lane="2" points="283" resultid="142" swimtime="00:00:44.62"><SPLITS/></RESULT><RESULT eventid="9" heatid="119" lane="6" points="366" resultid="901" swimtime="00:00:33.09"><SPLITS/></RESULT><RESULT eventid="11" heatid="164" lane="8" points="283" resultid="1242" swimtime="00:03:11.94"><SPLITS><SPLIT distance="50" swimtime="00:00:40.54"/><SPLIT distance="100" swimtime="00:01:30.58"/><SPLIT distance="150" swimtime="00:02:29.90"/></SPLITS></RESULT><RESULT eventid="31" heatid="338" lane="1" points="281" resultid="2515" swimtime="00:01:37.81"><SPLITS><SPLIT distance="50" swimtime="00:00:46.76"/></SPLITS></RESULT><RESULT eventid="35" heatid="376" lane="6" points="323" resultid="2803" swimtime="00:00:35.57"><SPLITS/></RESULT><RESULT eventid="39" heatid="435" lane="2" points="321" resultid="3243" swimtime="00:01:15.51"><SPLITS><SPLIT distance="50" swimtime="00:00:35.53"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="330" birthdate="2010-01-01" firstname="Sarah" gender="F" lastname="Kindseder" license="417858"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="45" lane="2" points="332" resultid="337" swimtime="00:05:41.13"><SPLITS><SPLIT distance="100" swimtime="00:01:19.46"/><SPLIT distance="200" swimtime="00:02:50.39"/><SPLIT distance="300" swimtime="00:04:15.53"/></SPLITS></RESULT><RESULT eventid="9" heatid="122" lane="8" points="352" resultid="927" swimtime="00:00:33.52"><SPLITS/></RESULT><RESULT eventid="13" heatid="201" lane="3" points="328" resultid="1522" swimtime="00:01:23.24"><SPLITS><SPLIT distance="50" swimtime="00:00:39.21"/></SPLITS></RESULT><RESULT eventid="27" heatid="269" lane="8" points="371" resultid="2002" swimtime="00:00:37.54"><SPLITS/></RESULT><RESULT eventid="31" heatid="336" lane="6" points="191" resultid="2504" swimtime="00:01:51.35"><SPLITS><SPLIT distance="50" swimtime="00:00:49.23"/></SPLITS></RESULT><RESULT eventid="35" heatid="372" lane="4" points="296" resultid="2770" swimtime="00:00:36.62"><SPLITS/></RESULT><RESULT eventid="39" heatid="440" lane="7" points="378" resultid="3287" swimtime="00:01:11.49"><SPLITS><SPLIT distance="50" swimtime="00:00:34.29"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="523" birthdate="2006-01-01" firstname="Vanessa" gender="F" lastname="Blaschke" license="387872"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="9" heatid="123" lane="2" points="394" resultid="929" swimtime="00:00:32.28"><SPLITS/></RESULT><RESULT eventid="13" heatid="207" lane="1" points="342" resultid="1568" swimtime="00:01:22.15"><SPLITS><SPLIT distance="50" swimtime="00:00:38.09"/></SPLITS></RESULT><RESULT eventid="27" heatid="271" lane="5" points="474" resultid="2014" swimtime="00:00:34.59"><SPLITS/></RESULT><RESULT eventid="35" heatid="378" lane="6" points="330" resultid="2817" swimtime="00:00:35.33"><SPLITS/></RESULT><RESULT eventid="39" heatid="443" lane="1" points="325" resultid="3305" swimtime="00:01:15.14"><SPLITS><SPLIT distance="50" swimtime="00:00:34.94"/></SPLITS></RESULT></RESULTS></ATHLETE></ATHLETES><RELAYS/></CLUB><CLUB code="4292" name="SC Prinz Eugen München" nation="GER" region="02" shortname="SCPE" type="CLUB"><CONTACT city="München" email="cheftrainer.schwimmen@scpe.de" fax="+49 89 625 7238" name="Mangafic, Elvir" phone="089 / 625 7238" street="Marianne-Plehn-Str. 23" zip="81825"/><OFFICIALS/><ATHLETES><ATHLETE athleteid="117" birthdate="2015-01-01" firstname="Marlene" gender="F" lastname="Berninger" license="471473"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="16" lane="1" points="248" resultid="117" swimtime="00:00:46.59"><SPLITS/></RESULT><RESULT eventid="7" heatid="86" lane="8" points="299" resultid="648" swimtime="00:03:27.57"><SPLITS><SPLIT distance="50" swimtime="00:00:48.24"/><SPLIT distance="100" swimtime="00:01:39.63"/><SPLIT distance="150" swimtime="00:02:35.06"/></SPLITS></RESULT><RESULT eventid="11" heatid="162" lane="8" points="262" resultid="1226" swimtime="00:03:16.86"><SPLITS><SPLIT distance="50" swimtime="00:00:47.49"/><SPLIT distance="100" swimtime="00:01:37.45"/><SPLIT distance="150" swimtime="00:02:31.50"/></SPLITS></RESULT><RESULT eventid="13" heatid="197" lane="1" points="194" resultid="1488" swimtime="00:01:39.15"><SPLITS><SPLIT distance="50" swimtime="00:00:47.59"/></SPLITS></RESULT><RESULT eventid="29" heatid="294" lane="1" points="231" resultid="2182" swimtime="00:03:04.09"><SPLITS><SPLIT distance="50" swimtime="00:00:40.67"/><SPLIT distance="100" swimtime="00:01:28.10"/><SPLIT distance="150" swimtime="00:02:18.10"/></SPLITS></RESULT><RESULT comment="12:31 Die Sportlerin hat nicht die vollständige Wettkampfstrecke absolviert" eventid="31" heatid="337" lane="5" resultid="2511" status="DSQ" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="125" birthdate="2013-01-01" firstname="Selma" gender="F" lastname="Schiermeier" license="492796"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="17" lane="1" resultid="125" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="7" heatid="86" lane="4" resultid="644" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="9" heatid="113" lane="7" resultid="855" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="159" birthdate="2008-01-01" firstname="Hanna" gender="F" lastname="Büttner" license="437861"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="21" lane="3" points="330" resultid="159" swimtime="00:00:42.37"><SPLITS/></RESULT><RESULT eventid="13" heatid="201" lane="5" points="258" resultid="1524" swimtime="00:01:30.19"><SPLITS><SPLIT distance="50" swimtime="00:00:43.10"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="170" birthdate="2007-01-01" firstname="Anna-Maria" gender="F" lastname="Kruse" license="388055"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="22" lane="8" points="295" resultid="170" swimtime="00:00:43.99"><SPLITS/></RESULT><RESULT eventid="5" heatid="67" lane="8" points="297" resultid="503" swimtime="00:01:23.11"><SPLITS><SPLIT distance="50" swimtime="00:00:37.53"/></SPLITS></RESULT><RESULT eventid="13" heatid="206" lane="7" points="343" resultid="1566" swimtime="00:01:22.04"><SPLITS><SPLIT distance="50" swimtime="00:00:39.48"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="219" birthdate="2014-01-01" firstname="Luca Mathias" gender="M" lastname="Kruse" license="451669"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="29" lane="7" points="127" resultid="219" swimtime="00:00:51.52"><SPLITS/></RESULT><RESULT eventid="10" heatid="137" lane="1" points="121" resultid="1029" swimtime="00:00:42.27"><SPLITS/></RESULT><RESULT eventid="14" heatid="212" lane="1" points="102" resultid="1605" swimtime="00:01:50.35"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="251" birthdate="2013-01-01" firstname="Francisko" gender="M" lastname="Linares Fernandez" license="461469"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="33" lane="7" points="204" resultid="251" swimtime="00:00:44.08"><SPLITS/></RESULT><RESULT eventid="8" heatid="98" lane="2" points="229" resultid="735" swimtime="00:03:25.64"><SPLITS><SPLIT distance="50" swimtime="00:00:45.01"/><SPLIT distance="100" swimtime="00:01:38.05"/><SPLIT distance="150" swimtime="00:02:31.85"/></SPLITS></RESULT><RESULT eventid="14" heatid="217" lane="3" points="182" resultid="1645" swimtime="00:01:31.00"><SPLITS><SPLIT distance="50" swimtime="00:00:44.78"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="255" birthdate="2013-01-01" firstname="Leon" gender="M" lastname="Starzynski" license="461470"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="34" lane="3" resultid="255" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="8" heatid="96" lane="2" resultid="719" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="10" heatid="141" lane="6" resultid="1064" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="14" heatid="218" lane="8" resultid="1658" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="260" birthdate="2012-01-01" firstname="Dmytro" gender="M" lastname="Pavlenko" license="460385"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="35" lane="2" points="201" resultid="260" swimtime="00:00:44.24"><SPLITS/></RESULT><RESULT eventid="12" heatid="183" lane="8" points="250" resultid="1388" swimtime="00:03:00.94"><SPLITS><SPLIT distance="50" swimtime="00:00:39.79"/><SPLIT distance="100" swimtime="00:01:25.92"/><SPLIT distance="150" swimtime="00:02:20.00"/></SPLITS></RESULT><RESULT eventid="14" heatid="219" lane="3" points="214" resultid="1661" swimtime="00:01:26.17"><SPLITS><SPLIT distance="50" swimtime="00:00:43.01"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="268" birthdate="2010-01-01" firstname="Noah" gender="M" lastname="Kaiser" license="463687"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="36" lane="2" points="305" resultid="268" swimtime="00:00:38.52"><SPLITS/></RESULT><RESULT eventid="8" heatid="99" lane="1" points="293" resultid="741" swimtime="00:03:09.45"><SPLITS><SPLIT distance="50" swimtime="00:00:43.89"/><SPLIT distance="100" swimtime="00:01:32.82"/><SPLIT distance="150" swimtime="00:02:21.03"/></SPLITS></RESULT><RESULT eventid="10" heatid="146" lane="2" points="311" resultid="1099" swimtime="00:00:30.85"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="277" birthdate="2009-01-01" firstname="Anir" gender="M" lastname="Bach-El Arif" license="466698"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="37" lane="3" points="309" resultid="277" swimtime="00:00:38.38"><SPLITS/></RESULT><RESULT eventid="10" heatid="148" lane="4" points="360" resultid="1117" swimtime="00:00:29.38"><SPLITS/></RESULT><RESULT eventid="32" heatid="353" lane="2" resultid="2628" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="36" heatid="395" lane="5" resultid="2946" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="40" heatid="468" lane="8" resultid="3505" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="283" birthdate="2008-01-01" firstname="Paul" gender="M" lastname="Rodionov" license="373312"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="38" lane="1" points="310" resultid="283" swimtime="00:00:38.33"><SPLITS/></RESULT><RESULT eventid="8" heatid="99" lane="3" points="296" resultid="743" swimtime="00:03:08.84"><SPLITS><SPLIT distance="50" swimtime="00:00:40.82"/><SPLIT distance="100" swimtime="00:01:29.25"/><SPLIT distance="150" swimtime="00:02:21.01"/></SPLITS></RESULT><RESULT eventid="10" heatid="152" lane="6" points="450" resultid="1151" swimtime="00:00:27.27"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="306" birthdate="2007-01-01" firstname="Maximilian" gender="M" lastname="Mühlbauer" license="390151"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="40" lane="8" points="534" resultid="306" swimtime="00:00:31.97"><SPLITS/></RESULT><RESULT eventid="6" heatid="79" lane="5" points="473" resultid="594" swimtime="00:01:03.43"><SPLITS><SPLIT distance="50" swimtime="00:00:28.40"/></SPLITS></RESULT><RESULT eventid="10" heatid="154" lane="7" points="490" resultid="1167" swimtime="00:00:26.52"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="358" birthdate="2009-01-01" firstname="Annabella" gender="F" lastname="E.C. Dullinger" license="454686"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="50" lane="2" points="372" resultid="376" swimtime="00:05:28.62"><SPLITS><SPLIT distance="100" swimtime="00:01:12.66"/><SPLIT distance="200" swimtime="00:02:34.68"/><SPLIT distance="300" swimtime="00:04:02.32"/></SPLITS></RESULT><RESULT eventid="29" heatid="303" lane="3" points="404" resultid="2255" swimtime="00:02:32.72"><SPLITS><SPLIT distance="50" swimtime="00:00:33.86"/><SPLIT distance="100" swimtime="00:01:12.94"/><SPLIT distance="150" swimtime="00:01:56.00"/></SPLITS></RESULT><RESULT eventid="39" heatid="444" lane="1" points="417" resultid="3313" swimtime="00:01:09.17"><SPLITS><SPLIT distance="50" swimtime="00:00:33.19"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="407" birthdate="2010-01-01" firstname="Kirill" gender="M" lastname="Lytschmann" license="413523"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="58" lane="2" points="314" resultid="435" swimtime="00:05:23.59"><SPLITS><SPLIT distance="100" swimtime="00:01:16.00"/><SPLIT distance="200" swimtime="00:02:40.28"/><SPLIT distance="300" swimtime="00:04:02.81"/></SPLITS></RESULT><RESULT eventid="8" heatid="99" lane="8" points="278" resultid="748" swimtime="00:03:12.80"><SPLITS><SPLIT distance="50" swimtime="00:00:45.04"/><SPLIT distance="100" swimtime="00:01:33.75"/><SPLIT distance="150" swimtime="00:02:24.63"/></SPLITS></RESULT><RESULT eventid="12" heatid="184" lane="2" points="299" resultid="1390" swimtime="00:02:50.48"><SPLITS><SPLIT distance="50" swimtime="00:00:37.81"/><SPLIT distance="100" swimtime="00:01:21.64"/><SPLIT distance="150" swimtime="00:02:12.42"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="412" birthdate="2013-01-01" firstname="David" gender="M" lastname="Rangelov" license="453834"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="59" lane="1" points="307" resultid="441" swimtime="00:05:25.93"><SPLITS><SPLIT distance="100" swimtime="00:01:14.44"/><SPLIT distance="200" swimtime="00:02:37.37"/><SPLIT distance="300" swimtime="00:04:03.28"/></SPLITS></RESULT><RESULT eventid="12" heatid="185" lane="2" points="310" resultid="1397" swimtime="00:02:48.32"><SPLITS><SPLIT distance="50" swimtime="00:00:36.01"/><SPLIT distance="100" swimtime="00:01:19.27"/><SPLIT distance="150" swimtime="00:02:11.20"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="460" birthdate="2010-01-01" firstname="Nila" gender="F" lastname="Schmidt-Hoensdorf" license="430267"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="5" heatid="70" lane="6" points="487" resultid="525" swimtime="00:01:10.48"><SPLITS><SPLIT distance="50" swimtime="00:00:32.07"/></SPLITS></RESULT><RESULT eventid="9" heatid="130" lane="5" points="551" resultid="987" swimtime="00:00:28.87"><SPLITS/></RESULT><RESULT eventid="33" heatid="360" lane="8" points="411" resultid="2682" swimtime="00:02:43.76"><SPLITS><SPLIT distance="50" swimtime="00:00:34.09"/><SPLIT distance="100" swimtime="00:01:13.14"/><SPLIT distance="150" swimtime="00:01:58.81"/></SPLITS></RESULT><RESULT eventid="35" heatid="382" lane="8" points="466" resultid="2851" swimtime="00:00:31.49"><SPLITS/></RESULT><RESULT eventid="39" heatid="449" lane="5" points="562" resultid="3354" swimtime="00:01:02.66"><SPLITS><SPLIT distance="50" swimtime="00:00:30.07"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="466" birthdate="2009-01-01" firstname="Mira" gender="F" lastname="Kolbmann" license="371264"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="5" heatid="71" lane="6" points="519" resultid="533" swimtime="00:01:09.03"><SPLITS><SPLIT distance="50" swimtime="00:00:31.45"/></SPLITS></RESULT><RESULT eventid="7" heatid="92" lane="4" points="635" resultid="692" swimtime="00:02:41.59"><SPLITS><SPLIT distance="50" swimtime="00:00:35.79"/><SPLIT distance="100" swimtime="00:01:17.09"/><SPLIT distance="150" swimtime="00:02:00.19"/></SPLITS></RESULT><RESULT eventid="11" heatid="174" lane="4" points="606" resultid="1318" swimtime="00:02:28.96"><SPLITS><SPLIT distance="50" swimtime="00:00:31.89"/><SPLIT distance="100" swimtime="00:01:11.46"/><SPLIT distance="150" swimtime="00:01:53.08"/></SPLITS></RESULT><RESULT eventid="13" heatid="209" lane="4" points="512" resultid="1586" swimtime="00:01:11.78"><SPLITS><SPLIT distance="50" swimtime="00:00:34.28"/></SPLITS></RESULT><RESULT eventid="31" heatid="344" lane="4" points="609" resultid="2566" swimtime="00:01:15.65"><SPLITS><SPLIT distance="50" swimtime="00:00:35.06"/></SPLITS></RESULT><RESULT eventid="33" heatid="360" lane="3" points="512" resultid="2677" swimtime="00:02:32.24"><SPLITS><SPLIT distance="50" swimtime="00:00:33.15"/><SPLIT distance="100" swimtime="00:01:11.21"/><SPLIT distance="150" swimtime="00:01:51.95"/></SPLITS></RESULT><RESULT eventid="37" heatid="412" lane="5" points="597" resultid="3075" swimtime="00:02:26.45"><SPLITS><SPLIT distance="100" swimtime="00:01:11.89"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="477" birthdate="2011-01-01" firstname="An-Simon" gender="M" lastname="Schmiegelt" license="467121"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="6" heatid="74" lane="5" points="166" resultid="555" swimtime="00:01:29.81"><SPLITS><SPLIT distance="50" swimtime="00:00:38.07"/></SPLITS></RESULT><RESULT eventid="10" heatid="147" lane="2" points="321" resultid="1107" swimtime="00:00:30.51"><SPLITS/></RESULT><RESULT eventid="14" heatid="222" lane="3" points="322" resultid="1684" swimtime="00:01:15.23"><SPLITS><SPLIT distance="50" swimtime="00:00:37.55"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="502" birthdate="2008-01-01" firstname="Leopold" gender="M" lastname="Becker" license="380655"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="6" heatid="80" lane="5" points="558" resultid="601" swimtime="00:01:00.04"><SPLITS><SPLIT distance="50" swimtime="00:00:28.41"/></SPLITS></RESULT><RESULT eventid="10" heatid="156" lane="2" points="537" resultid="1177" swimtime="00:00:25.71"><SPLITS/></RESULT><RESULT eventid="34" heatid="362" lane="4" points="561" resultid="2692" swimtime="00:02:13.77"><SPLITS><SPLIT distance="50" swimtime="00:00:28.88"/><SPLIT distance="100" swimtime="00:01:04.34"/><SPLIT distance="150" swimtime="00:01:40.01"/></SPLITS></RESULT><RESULT eventid="36" heatid="400" lane="4" points="590" resultid="2984" swimtime="00:00:26.55"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="558" birthdate="2008-01-01" firstname="Peter" gender="M" lastname="Rodionov" license="373313"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="10" heatid="155" lane="2" resultid="1170" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="12" heatid="188" lane="1" resultid="1420" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="14" heatid="223" lane="6" resultid="1695" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="562" birthdate="2011-01-01" firstname="Emma" gender="F" lastname="Vasilic" license="420144"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="11" heatid="174" lane="7" points="525" resultid="1321" swimtime="00:02:36.30"><SPLITS><SPLIT distance="50" swimtime="00:00:32.18"/><SPLIT distance="100" swimtime="00:01:11.82"/><SPLIT distance="150" swimtime="00:02:00.09"/></SPLITS></RESULT><RESULT eventid="13" heatid="209" lane="3" points="515" resultid="1585" swimtime="00:01:11.65"><SPLITS><SPLIT distance="50" swimtime="00:00:35.74"/></SPLITS></RESULT><RESULT eventid="27" heatid="272" lane="3" points="531" resultid="2020" swimtime="00:00:33.30"><SPLITS/></RESULT><RESULT eventid="29" heatid="306" lane="7" points="526" resultid="2281" swimtime="00:02:19.96"><SPLITS><SPLIT distance="50" swimtime="00:00:33.02"/><SPLIT distance="100" swimtime="00:01:08.72"/><SPLIT distance="150" swimtime="00:01:44.85"/></SPLITS></RESULT><RESULT eventid="37" heatid="412" lane="2" points="487" resultid="3072" swimtime="00:02:36.70"><SPLITS><SPLIT distance="100" swimtime="00:01:16.73"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="596" birthdate="2010-01-01" firstname="Maximilian" gender="M" lastname="Mansmann" license="394784"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="28" heatid="286" lane="2" points="420" resultid="2125" swimtime="00:00:31.65"><SPLITS/></RESULT><RESULT eventid="36" heatid="397" lane="2" points="455" resultid="2959" swimtime="00:00:28.94"><SPLITS/></RESULT><RESULT eventid="40" heatid="471" lane="7" points="417" resultid="3528" swimtime="00:01:02.70"><SPLITS><SPLIT distance="50" swimtime="00:00:29.23"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="597" birthdate="2008-01-01" firstname="Aleksej" gender="M" lastname="Brkic" license="419934"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="28" heatid="286" lane="7" points="399" resultid="2130" swimtime="00:00:32.19"><SPLITS/></RESULT><RESULT eventid="30" heatid="324" lane="2" points="439" resultid="2412" swimtime="00:02:14.17"><SPLITS><SPLIT distance="50" swimtime="00:00:29.19"/><SPLIT distance="100" swimtime="00:01:02.94"/><SPLIT distance="150" swimtime="00:01:38.05"/></SPLITS></RESULT><RESULT eventid="36" heatid="397" lane="7" points="452" resultid="2964" swimtime="00:00:29.00"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="606" birthdate="2008-01-01" firstname="Simon" gender="M" lastname="Metzger" license="444308"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="32" heatid="354" lane="2" points="297" resultid="2636" swimtime="00:01:25.19"><SPLITS><SPLIT distance="50" swimtime="00:00:40.38"/></SPLITS></RESULT><RESULT eventid="36" heatid="394" lane="1" points="290" resultid="2934" swimtime="00:00:33.61"><SPLITS/></RESULT><RESULT eventid="40" heatid="471" lane="6" points="384" resultid="3527" swimtime="00:01:04.46"><SPLITS><SPLIT distance="50" swimtime="00:00:30.23"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="607" birthdate="2008-01-01" firstname="Benedikt" gender="M" lastname="Weihe" license="449203"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="32" heatid="355" lane="6" points="409" resultid="2647" swimtime="00:01:16.62"><SPLITS><SPLIT distance="50" swimtime="00:00:36.47"/></SPLITS></RESULT><RESULT eventid="40" heatid="474" lane="7" points="531" resultid="3551" swimtime="00:00:57.86"><SPLITS><SPLIT distance="50" swimtime="00:00:27.86"/></SPLITS></RESULT></RESULTS></ATHLETE></ATHLETES><RELAYS><RELAY agemax="-1" agemin="-1" agetotalmax="17" agetotalmin="17" gender="F" name="1. Mannschaft" number="1"><ENTRIES/><RESULTS><RESULT eventid="43" heatid="482" lane="4" points="487" resultid="3598" swimtime="00:09:43.55"><SPLITS><SPLIT distance="50" swimtime="00:00:33.96"/><SPLIT distance="100" swimtime="00:01:14.58"/><SPLIT distance="150" swimtime="00:01:55.99"/><SPLIT distance="200" swimtime="00:02:38.54"/><SPLIT distance="250" swimtime="00:03:10.67"/><SPLIT distance="300" swimtime="00:03:46.45"/><SPLIT distance="350" swimtime="00:04:23.68"/><SPLIT distance="400" swimtime="00:05:00.59"/><SPLIT distance="450" swimtime="00:05:31.60"/><SPLIT distance="500" swimtime="00:06:09.44"/><SPLIT distance="550" swimtime="00:06:48.10"/><SPLIT distance="600" swimtime="00:07:25.53"/><SPLIT distance="650" swimtime="00:07:57.13"/><SPLIT distance="700" swimtime="00:08:33.01"/><SPLIT distance="750" swimtime="00:09:09.37"/></SPLITS><RELAYPOSITIONS><RELAYPOSITION athleteid="358" number="1"/><RELAYPOSITION athleteid="562" number="2"/><RELAYPOSITION athleteid="460" number="3"/><RELAYPOSITION athleteid="466" number="4"/></RELAYPOSITIONS></RESULT></RESULTS></RELAY></RELAYS></CLUB><CLUB code="PAZ" name="PLAVECKÁ AKADEMIE ZBUCH" nation="CZE" shortname="PAZ" type="CLUB"><CONTACT city="Plzen" country="CZE" email="vaclav.cermak@volny.cz" name="Cermák Václav" street="Krašovská 22" zip="32300"/><OFFICIALS/><ATHLETES><ATHLETE athleteid="144" birthdate="2010-01-01" firstname="Johanka" gender="F" lastname="Duchková" license="63450075"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="19" lane="4" points="376" resultid="144" swimtime="00:00:40.58"><SPLITS/></RESULT><RESULT eventid="7" heatid="89" lane="6" points="347" resultid="670" swimtime="00:03:17.55"><SPLITS><SPLIT distance="50" swimtime="00:00:46.14"/><SPLIT distance="100" swimtime="00:01:37.44"/><SPLIT distance="150" swimtime="00:02:28.92"/></SPLITS></RESULT><RESULT eventid="9" heatid="120" lane="4" points="385" resultid="907" swimtime="00:00:32.53"><SPLITS/></RESULT><RESULT eventid="17" heatid="230" lane="6" points="334" resultid="1737" swimtime="00:11:38.58"><SPLITS><SPLIT distance="100" swimtime="00:01:26.57"/><SPLIT distance="200" swimtime="00:02:56.71"/><SPLIT distance="300" swimtime="00:04:23.39"/><SPLIT distance="400" swimtime="00:05:50.10"/><SPLIT distance="500" swimtime="00:07:17.64"/><SPLIT distance="600" swimtime="00:08:45.91"/><SPLIT distance="700" swimtime="00:10:13.79"/></SPLITS></RESULT><RESULT eventid="29" heatid="299" lane="6" points="345" resultid="2227" swimtime="00:02:41.03"><SPLITS><SPLIT distance="50" swimtime="00:00:37.69"/><SPLIT distance="100" swimtime="00:01:19.18"/><SPLIT distance="150" swimtime="00:02:00.58"/></SPLITS></RESULT><RESULT eventid="31" heatid="340" lane="7" points="332" resultid="2537" swimtime="00:01:32.60"><SPLITS><SPLIT distance="50" swimtime="00:00:43.36"/></SPLITS></RESULT><RESULT eventid="35" heatid="371" lane="4" points="281" resultid="2762" swimtime="00:00:37.29"><SPLITS/></RESULT><RESULT eventid="39" heatid="439" lane="3" points="323" resultid="3276" swimtime="00:01:15.31"><SPLITS><SPLIT distance="50" swimtime="00:00:36.29"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="147" birthdate="2011-01-01" firstname="Barbora" gender="F" lastname="ŠKábová" license="63458611"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="19" lane="7" points="347" resultid="147" swimtime="00:00:41.66"><SPLITS/></RESULT><RESULT eventid="5" heatid="68" lane="4" points="400" resultid="507" swimtime="00:01:15.27"><SPLITS><SPLIT distance="50" swimtime="00:00:33.55"/></SPLITS></RESULT><RESULT eventid="9" heatid="128" lane="3" points="444" resultid="969" swimtime="00:00:31.01"><SPLITS/></RESULT><RESULT eventid="11" heatid="170" lane="4" points="446" resultid="1286" swimtime="00:02:45.03"><SPLITS><SPLIT distance="50" swimtime="00:00:35.65"/><SPLIT distance="100" swimtime="00:01:20.31"/><SPLIT distance="150" swimtime="00:02:08.31"/></SPLITS></RESULT><RESULT eventid="13" heatid="204" lane="8" points="376" resultid="1551" swimtime="00:01:19.55"><SPLITS><SPLIT distance="50" swimtime="00:00:39.10"/></SPLITS></RESULT><RESULT eventid="29" heatid="304" lane="6" points="466" resultid="2266" swimtime="00:02:25.63"><SPLITS><SPLIT distance="50" swimtime="00:00:32.97"/><SPLIT distance="100" swimtime="00:01:09.67"/><SPLIT distance="150" swimtime="00:01:47.51"/></SPLITS></RESULT><RESULT eventid="33" heatid="359" lane="5" points="319" resultid="2671" swimtime="00:02:58.25"><SPLITS><SPLIT distance="50" swimtime="00:00:37.07"/><SPLIT distance="100" swimtime="00:01:20.64"/><SPLIT distance="150" swimtime="00:02:09.01"/></SPLITS></RESULT><RESULT eventid="35" heatid="375" lane="5" points="393" resultid="2794" swimtime="00:00:33.33"><SPLITS/></RESULT><RESULT eventid="41" heatid="478" lane="8" points="400" resultid="3577" swimtime="00:06:01.36"><SPLITS><SPLIT distance="50" swimtime="00:00:38.50"/><SPLIT distance="100" swimtime="00:01:25.54"/><SPLIT distance="150" swimtime="00:02:13.10"/><SPLIT distance="200" swimtime="00:02:58.19"/><SPLIT distance="250" swimtime="00:03:49.61"/><SPLIT distance="300" swimtime="00:04:41.07"/><SPLIT distance="350" swimtime="00:05:21.55"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="291" birthdate="2010-01-01" firstname="Vilém" gender="M" lastname="Hanzel" license="52095000"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="39" lane="1" points="372" resultid="291" swimtime="00:00:36.08"><SPLITS/></RESULT><RESULT eventid="6" heatid="79" lane="7" points="489" resultid="596" swimtime="00:01:02.74"><SPLITS><SPLIT distance="50" swimtime="00:00:28.95"/></SPLITS></RESULT><RESULT eventid="10" heatid="154" lane="4" points="469" resultid="1165" swimtime="00:00:26.91"><SPLITS/></RESULT><RESULT eventid="12" heatid="188" lane="3" points="415" resultid="1422" swimtime="00:02:32.80"><SPLITS><SPLIT distance="50" swimtime="00:00:30.67"/><SPLIT distance="100" swimtime="00:01:12.01"/><SPLIT distance="150" swimtime="00:01:57.72"/></SPLITS></RESULT><RESULT eventid="32" heatid="355" lane="5" points="397" resultid="2646" swimtime="00:01:17.36"><SPLITS><SPLIT distance="50" swimtime="00:00:35.56"/></SPLITS></RESULT><RESULT eventid="34" heatid="362" lane="2" points="325" resultid="2690" swimtime="00:02:40.44"><SPLITS><SPLIT distance="50" swimtime="00:00:32.46"/><SPLIT distance="100" swimtime="00:01:10.91"/><SPLIT distance="150" swimtime="00:01:54.60"/></SPLITS></RESULT><RESULT eventid="36" heatid="398" lane="5" points="501" resultid="2970" swimtime="00:00:28.03"><SPLITS/></RESULT><RESULT eventid="40" heatid="473" lane="4" points="514" resultid="3540" swimtime="00:00:58.48"><SPLITS><SPLIT distance="50" swimtime="00:00:27.47"/></SPLITS></RESULT><RESULT eventid="42" heatid="480" lane="6" points="320" resultid="3589" swimtime="00:05:56.27"><SPLITS><SPLIT distance="50" swimtime="00:00:36.86"/><SPLIT distance="100" swimtime="00:01:20.42"/><SPLIT distance="150" swimtime="00:02:08.54"/><SPLIT distance="200" swimtime="00:02:55.55"/><SPLIT distance="250" swimtime="00:03:47.03"/><SPLIT distance="300" swimtime="00:04:37.88"/><SPLIT distance="350" swimtime="00:05:17.32"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="356" birthdate="2009-01-01" firstname="Karolína" gender="F" lastname="Šmídovcová" license="54424000"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="49" lane="8" points="342" resultid="374" swimtime="00:05:37.93"><SPLITS><SPLIT distance="100" swimtime="00:01:12.78"/><SPLIT distance="200" swimtime="00:02:38.56"/><SPLIT distance="300" swimtime="00:04:08.53"/></SPLITS></RESULT><RESULT eventid="9" heatid="124" lane="5" points="419" resultid="940" swimtime="00:00:31.63"><SPLITS/></RESULT><RESULT eventid="13" heatid="206" lane="6" points="387" resultid="1565" swimtime="00:01:18.77"><SPLITS><SPLIT distance="50" swimtime="00:00:38.29"/></SPLITS></RESULT><RESULT eventid="17" heatid="231" lane="7" points="354" resultid="1746" swimtime="00:11:24.70"><SPLITS><SPLIT distance="100" swimtime="00:01:15.26"/><SPLIT distance="200" swimtime="00:02:38.97"/><SPLIT distance="300" swimtime="00:04:05.05"/><SPLIT distance="400" swimtime="00:05:32.52"/><SPLIT distance="500" swimtime="00:07:00.37"/><SPLIT distance="600" swimtime="00:08:29.08"/><SPLIT distance="700" swimtime="00:09:58.60"/></SPLITS></RESULT><RESULT eventid="27" heatid="268" lane="5" points="397" resultid="1992" swimtime="00:00:36.69"><SPLITS/></RESULT><RESULT eventid="29" heatid="302" lane="3" points="369" resultid="2247" swimtime="00:02:37.49"><SPLITS><SPLIT distance="50" swimtime="00:00:34.94"/><SPLIT distance="100" swimtime="00:01:13.98"/><SPLIT distance="150" swimtime="00:01:56.07"/></SPLITS></RESULT><RESULT eventid="35" heatid="373" lane="5" points="336" resultid="2779" swimtime="00:00:35.11"><SPLITS/></RESULT><RESULT eventid="37" heatid="409" lane="6" points="345" resultid="3052" swimtime="00:02:55.80"><SPLITS><SPLIT distance="50" swimtime="00:00:38.92"/><SPLIT distance="100" swimtime="00:01:23.24"/><SPLIT distance="150" swimtime="00:02:08.68"/></SPLITS></RESULT><RESULT eventid="39" heatid="444" lane="5" points="396" resultid="3317" swimtime="00:01:10.38"><SPLITS><SPLIT distance="50" swimtime="00:00:33.01"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="424" birthdate="2009-01-01" firstname="Matej" gender="M" lastname="Flaks" license="49613000"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="60" lane="6" points="452" resultid="453" swimtime="00:04:46.66"><SPLITS><SPLIT distance="100" swimtime="00:01:07.82"/><SPLIT distance="200" swimtime="00:02:23.03"/><SPLIT distance="300" swimtime="00:03:38.00"/></SPLITS></RESULT><RESULT eventid="10" heatid="157" lane="4" points="614" resultid="1187" swimtime="00:00:24.59"><SPLITS/></RESULT><RESULT eventid="14" heatid="225" lane="5" points="584" resultid="1708" swimtime="00:01:01.70"><SPLITS><SPLIT distance="50" swimtime="00:00:29.99"/></SPLITS></RESULT><RESULT eventid="28" heatid="287" lane="5" points="594" resultid="2136" swimtime="00:00:28.20"><SPLITS/></RESULT><RESULT eventid="30" heatid="324" lane="5" points="424" resultid="2415" swimtime="00:02:15.71"><SPLITS><SPLIT distance="50" swimtime="00:00:28.91"/><SPLIT distance="100" swimtime="00:01:02.57"/><SPLIT distance="150" swimtime="00:01:39.75"/></SPLITS></RESULT><RESULT eventid="36" heatid="399" lane="6" points="532" resultid="2979" swimtime="00:00:27.47"><SPLITS/></RESULT><RESULT eventid="38" heatid="419" lane="5" points="410" resultid="3123" swimtime="00:02:30.62"><SPLITS><SPLIT distance="50" swimtime="00:00:33.55"/><SPLIT distance="100" swimtime="00:01:11.08"/><SPLIT distance="150" swimtime="00:01:52.39"/></SPLITS></RESULT><RESULT eventid="40" heatid="475" lane="6" points="498" resultid="3557" swimtime="00:00:59.08"><SPLITS><SPLIT distance="50" swimtime="00:00:27.62"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="427" birthdate="2009-01-01" firstname="Marek" gender="M" lastname="Šmídovec" license="54425000"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="61" lane="1" points="443" resultid="456" swimtime="00:04:48.50"><SPLITS><SPLIT distance="100" swimtime="00:01:02.74"/><SPLIT distance="200" swimtime="00:02:15.28"/><SPLIT distance="300" swimtime="00:03:32.18"/></SPLITS></RESULT><RESULT eventid="6" heatid="79" lane="4" points="454" resultid="593" swimtime="00:01:04.30"><SPLITS><SPLIT distance="50" swimtime="00:00:28.76"/></SPLITS></RESULT><RESULT eventid="10" heatid="156" lane="7" points="517" resultid="1182" swimtime="00:00:26.04"><SPLITS/></RESULT><RESULT eventid="30" heatid="324" lane="6" points="535" resultid="2416" swimtime="00:02:05.60"><SPLITS><SPLIT distance="50" swimtime="00:00:28.11"/><SPLIT distance="100" swimtime="00:00:59.35"/><SPLIT distance="150" swimtime="00:01:32.27"/></SPLITS></RESULT><RESULT eventid="34" heatid="362" lane="8" points="278" resultid="2695" swimtime="00:02:49.02"><SPLITS><SPLIT distance="50" swimtime="00:00:34.20"/><SPLIT distance="100" swimtime="00:01:16.08"/><SPLIT distance="150" swimtime="00:02:04.38"/></SPLITS></RESULT><RESULT eventid="36" heatid="399" lane="2" points="482" resultid="2975" swimtime="00:00:28.39"><SPLITS/></RESULT><RESULT eventid="40" heatid="474" lane="3" points="532" resultid="3547" swimtime="00:00:57.80"><SPLITS><SPLIT distance="50" swimtime="00:00:27.38"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="434" birthdate="2007-01-01" firstname="Petr" gender="M" lastname="Hajšman" license="54413000"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="62" lane="2" points="493" resultid="463" swimtime="00:04:38.43"><SPLITS><SPLIT distance="100" swimtime="00:01:00.28"/><SPLIT distance="200" swimtime="00:02:12.59"/><SPLIT distance="300" swimtime="00:03:26.58"/></SPLITS></RESULT><RESULT eventid="6" heatid="80" lane="1" points="440" resultid="598" swimtime="00:01:05.00"><SPLITS><SPLIT distance="50" swimtime="00:00:30.44"/></SPLITS></RESULT><RESULT eventid="10" heatid="157" lane="6" points="529" resultid="1189" swimtime="00:00:25.85"><SPLITS/></RESULT><RESULT eventid="30" heatid="325" lane="2" points="504" resultid="2420" swimtime="00:02:08.13"><SPLITS><SPLIT distance="50" swimtime="00:00:27.65"/><SPLIT distance="100" swimtime="00:01:00.17"/><SPLIT distance="150" swimtime="00:01:34.70"/></SPLITS></RESULT><RESULT eventid="36" heatid="399" lane="5" points="511" resultid="2978" swimtime="00:00:27.84"><SPLITS/></RESULT><RESULT eventid="40" heatid="475" lane="3" points="548" resultid="3554" swimtime="00:00:57.25"><SPLITS><SPLIT distance="50" swimtime="00:00:27.03"/></SPLITS></RESULT><RESULT eventid="42" heatid="481" lane="6" points="386" resultid="3595" swimtime="00:05:34.82"><SPLITS><SPLIT distance="50" swimtime="00:00:33.03"/><SPLIT distance="100" swimtime="00:01:14.44"/><SPLIT distance="150" swimtime="00:02:03.39"/><SPLIT distance="200" swimtime="00:02:47.46"/><SPLIT distance="250" swimtime="00:03:32.86"/><SPLIT distance="300" swimtime="00:04:19.66"/><SPLIT distance="350" swimtime="00:04:57.22"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="436" birthdate="2010-01-01" firstname="Adam" gender="M" lastname="Potucek" license="53461000"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="62" lane="6" points="525" resultid="466" swimtime="00:04:32.71"><SPLITS><SPLIT distance="100" swimtime="00:01:02.03"/><SPLIT distance="200" swimtime="00:02:11.75"/><SPLIT distance="300" swimtime="00:03:22.65"/></SPLITS></RESULT><RESULT eventid="6" heatid="79" lane="3" points="458" resultid="592" swimtime="00:01:04.15"><SPLITS><SPLIT distance="50" swimtime="00:00:29.52"/></SPLITS></RESULT><RESULT eventid="12" heatid="189" lane="6" points="491" resultid="1432" swimtime="00:02:24.50"><SPLITS><SPLIT distance="50" swimtime="00:00:28.75"/><SPLIT distance="100" swimtime="00:01:06.48"/><SPLIT distance="150" swimtime="00:01:52.13"/></SPLITS></RESULT><RESULT eventid="14" heatid="224" lane="8" points="376" resultid="1704" swimtime="00:01:11.48"><SPLITS><SPLIT distance="50" swimtime="00:00:34.87"/></SPLITS></RESULT><RESULT eventid="16" heatid="229" lane="5" points="500" resultid="1729" swimtime="00:18:17.19"><SPLITS><SPLIT distance="100" swimtime="00:01:05.63"/><SPLIT distance="200" swimtime="00:02:16.36"/><SPLIT distance="300" swimtime="00:03:27.34"/><SPLIT distance="400" swimtime="00:04:38.57"/><SPLIT distance="500" swimtime="00:05:50.56"/><SPLIT distance="600" swimtime="00:07:04.88"/><SPLIT distance="700" swimtime="00:08:19.14"/><SPLIT distance="800" swimtime="00:09:33.84"/><SPLIT distance="900" swimtime="00:10:48.62"/><SPLIT distance="1000" swimtime="00:12:03.95"/><SPLIT distance="1100" swimtime="00:13:19.08"/><SPLIT distance="1200" swimtime="00:14:34.47"/><SPLIT distance="1300" swimtime="00:15:49.61"/><SPLIT distance="1400" swimtime="00:17:03.85"/></SPLITS></RESULT><RESULT eventid="30" heatid="323" lane="4" points="493" resultid="2406" swimtime="00:02:09.09"><SPLITS><SPLIT distance="50" swimtime="00:00:28.44"/><SPLIT distance="100" swimtime="00:01:01.37"/><SPLIT distance="150" swimtime="00:01:35.57"/></SPLITS></RESULT><RESULT eventid="34" heatid="362" lane="6" points="299" resultid="2694" swimtime="00:02:44.83"><SPLITS><SPLIT distance="50" swimtime="00:00:31.73"/><SPLIT distance="100" swimtime="00:01:16.70"/><SPLIT distance="150" swimtime="00:02:03.83"/></SPLITS></RESULT><RESULT eventid="36" heatid="397" lane="4" points="464" resultid="2961" swimtime="00:00:28.75"><SPLITS/></RESULT><RESULT eventid="42" heatid="481" lane="3" points="460" resultid="3593" swimtime="00:05:15.75"><SPLITS><SPLIT distance="50" swimtime="00:00:30.11"/><SPLIT distance="100" swimtime="00:01:07.70"/><SPLIT distance="150" swimtime="00:01:50.81"/><SPLIT distance="200" swimtime="00:02:30.49"/><SPLIT distance="250" swimtime="00:03:18.17"/><SPLIT distance="300" swimtime="00:04:06.32"/><SPLIT distance="350" swimtime="00:04:41.54"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="444" birthdate="2012-01-01" firstname="Katerina" gender="F" lastname="Rašková" license="63440533"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="5" heatid="65" lane="2" points="198" resultid="482" swimtime="00:01:35.11"><SPLITS><SPLIT distance="50" swimtime="00:00:40.77"/></SPLITS></RESULT><RESULT eventid="9" heatid="118" lane="1" points="288" resultid="888" swimtime="00:00:35.81"><SPLITS/></RESULT><RESULT eventid="13" heatid="203" lane="6" points="298" resultid="1541" swimtime="00:01:26.01"><SPLITS><SPLIT distance="50" swimtime="00:00:41.26"/></SPLITS></RESULT><RESULT eventid="17" heatid="230" lane="2" points="308" resultid="1733" swimtime="00:11:57.49"><SPLITS><SPLIT distance="100" swimtime="00:01:21.51"/><SPLIT distance="200" swimtime="00:02:53.96"/><SPLIT distance="300" swimtime="00:04:26.03"/><SPLIT distance="400" swimtime="00:05:58.41"/><SPLIT distance="500" swimtime="00:07:29.65"/><SPLIT distance="600" swimtime="00:09:01.80"/><SPLIT distance="700" swimtime="00:10:32.61"/></SPLITS></RESULT><RESULT eventid="27" heatid="264" lane="6" points="300" resultid="1961" swimtime="00:00:40.27"><SPLITS/></RESULT><RESULT eventid="29" heatid="298" lane="3" points="308" resultid="2216" swimtime="00:02:47.16"><SPLITS><SPLIT distance="50" swimtime="00:00:37.35"/><SPLIT distance="100" swimtime="00:01:20.16"/><SPLIT distance="150" swimtime="00:02:06.51"/></SPLITS></RESULT><RESULT eventid="35" heatid="371" lane="1" points="213" resultid="2759" swimtime="00:00:40.88"><SPLITS/></RESULT><RESULT eventid="37" heatid="406" lane="5" points="309" resultid="3027" swimtime="00:03:02.38"><SPLITS><SPLIT distance="50" swimtime="00:00:42.32"/><SPLIT distance="100" swimtime="00:01:29.85"/><SPLIT distance="150" swimtime="00:02:17.93"/></SPLITS></RESULT><RESULT eventid="39" heatid="435" lane="5" points="282" resultid="3246" swimtime="00:01:18.83"><SPLITS><SPLIT distance="50" swimtime="00:00:37.15"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="504" birthdate="2010-01-01" firstname="Alexandr" gender="M" lastname="Beran" license="51975000"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="6" heatid="80" lane="7" points="506" resultid="603" swimtime="00:01:02.04"><SPLITS><SPLIT distance="50" swimtime="00:00:28.99"/></SPLITS></RESULT><RESULT eventid="10" heatid="157" lane="5" points="571" resultid="1188" swimtime="00:00:25.20"><SPLITS/></RESULT><RESULT eventid="30" heatid="325" lane="5" points="547" resultid="2422" swimtime="00:02:04.66"><SPLITS><SPLIT distance="50" swimtime="00:00:27.96"/><SPLIT distance="100" swimtime="00:00:59.28"/><SPLIT distance="150" swimtime="00:01:32.29"/></SPLITS></RESULT><RESULT eventid="36" heatid="400" lane="3" points="547" resultid="2983" swimtime="00:00:27.23"><SPLITS/></RESULT><RESULT eventid="40" heatid="475" lane="4" points="590" resultid="3555" swimtime="00:00:55.87"><SPLITS><SPLIT distance="50" swimtime="00:00:26.60"/></SPLITS></RESULT><RESULT eventid="42" heatid="480" lane="4" points="414" resultid="3588" swimtime="00:05:26.92"><SPLITS><SPLIT distance="50" swimtime="00:00:30.69"/><SPLIT distance="100" swimtime="00:01:10.51"/><SPLIT distance="150" swimtime="00:01:53.39"/><SPLIT distance="200" swimtime="00:02:36.59"/><SPLIT distance="250" swimtime="00:03:24.58"/><SPLIT distance="300" swimtime="00:04:15.88"/><SPLIT distance="350" swimtime="00:04:50.70"/></SPLITS></RESULT></RESULTS></ATHLETE></ATHLETES><RELAYS/></CLUB><CLUB code="6628" name="TSV Indersdorf" nation="GER" region="02" shortname="Indersdo" type="CLUB"><CONTACT city="Markt Indersdorf" country="GER" email="meldungen@indersdorfer-haie.de" name="Fett, Claudius-Franz" phone="08136 99214" street="Arnbacher Str 1" zip="85229"/><OFFICIALS/><ATHLETES><ATHLETE athleteid="161" birthdate="2011-01-01" firstname="Magdalena" gender="F" lastname="Kiefl" license="424453"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="21" lane="6" points="449" resultid="161" swimtime="00:00:38.24"><SPLITS/></RESULT><RESULT eventid="9" heatid="128" lane="1" points="478" resultid="967" swimtime="00:00:30.26"><SPLITS/></RESULT><RESULT eventid="13" heatid="204" lane="4" points="415" resultid="1547" swimtime="00:01:16.97"><SPLITS><SPLIT distance="50" swimtime="00:00:37.00"/></SPLITS></RESULT><RESULT eventid="27" heatid="266" lane="1" points="414" resultid="1972" swimtime="00:00:36.18"><SPLITS/></RESULT><RESULT eventid="37" heatid="409" lane="2" points="413" resultid="3048" swimtime="00:02:45.51"><SPLITS><SPLIT distance="50" swimtime="00:00:38.91"/><SPLIT distance="100" swimtime="00:01:21.59"/><SPLIT distance="150" swimtime="00:02:04.68"/></SPLITS></RESULT><RESULT eventid="39" heatid="445" lane="4" points="503" resultid="3324" swimtime="00:01:05.02"><SPLITS><SPLIT distance="50" swimtime="00:00:30.89"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="327" birthdate="2011-01-01" firstname="Emiliana" gender="F" lastname="Meretta Montoya" license="424456"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="44" lane="6" points="300" resultid="333" swimtime="00:05:53.00"><SPLITS><SPLIT distance="100" swimtime="00:01:23.25"/><SPLIT distance="200" swimtime="00:02:54.23"/><SPLIT distance="300" swimtime="00:04:26.06"/></SPLITS></RESULT><RESULT eventid="9" heatid="114" lane="3" points="338" resultid="859" swimtime="00:00:33.98"><SPLITS/></RESULT><RESULT eventid="13" heatid="201" lane="2" points="240" resultid="1521" swimtime="00:01:32.44"><SPLITS><SPLIT distance="50" swimtime="00:00:45.02"/></SPLITS></RESULT><RESULT eventid="15" heatid="226" lane="4" points="266" resultid="1715" swimtime="00:23:50.67"><SPLITS><SPLIT distance="100" swimtime="00:01:23.56"/><SPLIT distance="200" swimtime="00:02:57.99"/><SPLIT distance="300" swimtime="00:04:31.62"/><SPLIT distance="400" swimtime="00:06:07.16"/><SPLIT distance="500" swimtime="00:07:41.47"/><SPLIT distance="600" swimtime="00:09:19.01"/><SPLIT distance="700" swimtime="00:10:56.65"/><SPLIT distance="800" swimtime="00:12:33.48"/><SPLIT distance="900" swimtime="00:14:10.20"/><SPLIT distance="1000" swimtime="00:15:48.51"/><SPLIT distance="1100" swimtime="00:17:28.10"/><SPLIT distance="1200" swimtime="00:19:04.88"/><SPLIT distance="1300" swimtime="00:20:44.39"/><SPLIT distance="1400" swimtime="00:22:22.02"/></SPLITS></RESULT><RESULT eventid="27" heatid="263" lane="1" points="239" resultid="1948" swimtime="00:00:43.43"><SPLITS/></RESULT><RESULT eventid="35" heatid="371" lane="6" points="208" resultid="2764" swimtime="00:00:41.23"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="337" birthdate="2007-01-01" firstname="Paula" gender="F" lastname="Renhof" license="398238"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="46" lane="4" points="305" resultid="347" swimtime="00:05:51.01"><SPLITS><SPLIT distance="100" swimtime="00:01:21.05"/><SPLIT distance="200" swimtime="00:02:49.51"/><SPLIT distance="300" swimtime="00:04:20.75"/></SPLITS></RESULT><RESULT eventid="11" heatid="164" lane="7" points="265" resultid="1241" swimtime="00:03:16.11"><SPLITS><SPLIT distance="50" swimtime="00:00:42.39"/><SPLIT distance="100" swimtime="00:01:30.14"/><SPLIT distance="150" swimtime="00:02:32.17"/></SPLITS></RESULT><RESULT eventid="13" heatid="201" lane="7" points="260" resultid="1526" swimtime="00:01:30.00"><SPLITS><SPLIT distance="50" swimtime="00:00:43.51"/></SPLITS></RESULT><RESULT eventid="15" heatid="226" lane="1" points="283" resultid="1712" swimtime="00:23:21.42"><SPLITS><SPLIT distance="100" swimtime="00:01:24.08"/><SPLIT distance="200" swimtime="00:02:56.86"/><SPLIT distance="300" swimtime="00:04:29.92"/><SPLIT distance="400" swimtime="00:06:03.18"/><SPLIT distance="500" swimtime="00:07:36.41"/><SPLIT distance="600" swimtime="00:09:10.12"/><SPLIT distance="700" swimtime="00:10:43.89"/><SPLIT distance="800" swimtime="00:12:18.86"/><SPLIT distance="900" swimtime="00:13:53.21"/><SPLIT distance="1000" swimtime="00:15:28.18"/><SPLIT distance="1100" swimtime="00:17:02.90"/><SPLIT distance="1200" swimtime="00:18:38.04"/><SPLIT distance="1300" swimtime="00:20:13.00"/><SPLIT distance="1400" swimtime="00:21:48.02"/></SPLITS></RESULT><RESULT eventid="31" heatid="335" lane="3" points="209" resultid="2493" swimtime="00:01:47.97"><SPLITS><SPLIT distance="50" swimtime="00:00:52.29"/></SPLITS></RESULT><RESULT eventid="37" heatid="407" lane="7" points="290" resultid="3037" swimtime="00:03:06.34"><SPLITS><SPLIT distance="50" swimtime="00:00:43.39"/><SPLIT distance="100" swimtime="00:01:30.87"/><SPLIT distance="150" swimtime="00:02:19.07"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="442" birthdate="2012-01-01" firstname="Luisa" gender="F" lastname="Zangerle" license="437814"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="5" heatid="64" lane="6" points="278" resultid="478" swimtime="00:01:24.92"><SPLITS><SPLIT distance="50" swimtime="00:00:37.68"/></SPLITS></RESULT><RESULT eventid="13" heatid="201" lane="4" points="328" resultid="1523" swimtime="00:01:23.30"><SPLITS><SPLIT distance="50" swimtime="00:00:39.81"/></SPLITS></RESULT><RESULT eventid="27" heatid="267" lane="7" points="355" resultid="1986" swimtime="00:00:38.08"><SPLITS/></RESULT><RESULT eventid="29" heatid="297" lane="1" points="280" resultid="2206" swimtime="00:02:52.57"><SPLITS><SPLIT distance="50" swimtime="00:00:38.15"/><SPLIT distance="100" swimtime="00:01:21.87"/><SPLIT distance="150" swimtime="00:02:09.55"/></SPLITS></RESULT><RESULT eventid="35" heatid="373" lane="6" points="285" resultid="2780" swimtime="00:00:37.10"><SPLITS/></RESULT><RESULT eventid="37" heatid="406" lane="1" points="313" resultid="3023" swimtime="00:03:01.52"><SPLITS><SPLIT distance="50" swimtime="00:00:42.44"/><SPLIT distance="100" swimtime="00:01:29.04"/><SPLIT distance="150" swimtime="00:02:17.07"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="482" birthdate="2010-01-01" firstname="Felix" gender="M" lastname="Kannegießer" license="417940"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="6" heatid="75" lane="5" points="217" resultid="563" swimtime="00:01:22.28"><SPLITS><SPLIT distance="50" swimtime="00:00:34.89"/></SPLITS></RESULT><RESULT eventid="10" heatid="145" lane="2" points="351" resultid="1091" swimtime="00:00:29.63"><SPLITS/></RESULT><RESULT eventid="12" heatid="182" lane="1" points="266" resultid="1374" swimtime="00:02:57.08"><SPLITS><SPLIT distance="50" swimtime="00:00:38.68"/><SPLIT distance="100" swimtime="00:01:25.19"/><SPLIT distance="150" swimtime="00:02:17.36"/></SPLITS></RESULT><RESULT eventid="16" heatid="228" lane="8" points="340" resultid="1725" swimtime="00:20:46.95"><SPLITS><SPLIT distance="100" swimtime="00:01:13.05"/><SPLIT distance="200" swimtime="00:02:34.28"/><SPLIT distance="300" swimtime="00:03:57.49"/><SPLIT distance="400" swimtime="00:05:21.76"/><SPLIT distance="500" swimtime="00:06:46.81"/><SPLIT distance="600" swimtime="00:08:11.63"/><SPLIT distance="700" swimtime="00:09:35.34"/><SPLIT distance="800" swimtime="00:10:58.29"/><SPLIT distance="900" swimtime="00:12:21.98"/><SPLIT distance="1000" swimtime="00:13:44.68"/><SPLIT distance="1100" swimtime="00:15:07.86"/><SPLIT distance="1200" swimtime="00:16:31.06"/><SPLIT distance="1300" swimtime="00:17:57.16"/><SPLIT distance="1400" swimtime="00:19:23.28"/></SPLITS></RESULT><RESULT eventid="28" heatid="284" lane="7" resultid="2114" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="30" heatid="319" lane="2" resultid="2375" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="487" birthdate="2008-01-01" firstname="Ludwig" gender="M" lastname="Kost" license="385105"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="6" heatid="76" lane="7" points="308" resultid="573" swimtime="00:01:13.18"><SPLITS><SPLIT distance="50" swimtime="00:00:30.63"/></SPLITS></RESULT><RESULT eventid="10" heatid="157" lane="2" points="580" resultid="1185" swimtime="00:00:25.06"><SPLITS/></RESULT><RESULT eventid="14" heatid="223" lane="1" points="370" resultid="1690" swimtime="00:01:11.86"><SPLITS><SPLIT distance="50" swimtime="00:00:35.09"/></SPLITS></RESULT><RESULT eventid="16" heatid="229" lane="4" points="299" resultid="1728" swimtime="00:21:41.85"><SPLITS><SPLIT distance="100" swimtime="00:01:09.76"/><SPLIT distance="200" swimtime="00:02:31.75"/><SPLIT distance="300" swimtime="00:03:58.44"/><SPLIT distance="400" swimtime="00:05:27.91"/><SPLIT distance="500" swimtime="00:06:57.51"/><SPLIT distance="600" swimtime="00:08:28.12"/><SPLIT distance="700" swimtime="00:09:57.28"/><SPLIT distance="800" swimtime="00:11:27.64"/><SPLIT distance="900" swimtime="00:12:56.91"/><SPLIT distance="1000" swimtime="00:14:26.23"/><SPLIT distance="1100" swimtime="00:15:54.55"/><SPLIT distance="1200" swimtime="00:17:23.15"/><SPLIT distance="1300" swimtime="00:18:51.97"/><SPLIT distance="1400" swimtime="00:20:20.37"/></SPLITS></RESULT><RESULT eventid="36" heatid="397" lane="5" points="463" resultid="2962" swimtime="00:00:28.78"><SPLITS/></RESULT><RESULT eventid="40" heatid="473" lane="2" points="561" resultid="3538" swimtime="00:00:56.81"><SPLITS><SPLIT distance="50" swimtime="00:00:26.58"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="560" birthdate="2014-01-01" firstname="Valeria" gender="F" lastname="Meretta Montoya" license="472925"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="11" heatid="159" lane="4" points="175" resultid="1199" swimtime="00:03:45.07"><SPLITS><SPLIT distance="50" swimtime="00:00:53.52"/><SPLIT distance="100" swimtime="00:01:51.52"/><SPLIT distance="150" swimtime="00:02:54.16"/></SPLITS></RESULT><RESULT eventid="23" heatid="243" lane="6" resultid="1812" swimtime="00:00:57.03"><SPLITS/></RESULT><RESULT eventid="25" heatid="249" lane="7" resultid="1851" swimtime="00:01:04.57"><SPLITS/></RESULT><RESULT eventid="29" heatid="293" lane="4" points="186" resultid="2177" swimtime="00:03:17.77"><SPLITS><SPLIT distance="50" swimtime="00:00:42.79"/><SPLIT distance="100" swimtime="00:01:34.64"/><SPLIT distance="150" swimtime="00:02:29.69"/></SPLITS></RESULT><RESULT eventid="31" heatid="332" lane="3" points="183" resultid="2469" swimtime="00:01:52.83"><SPLITS><SPLIT distance="50" swimtime="00:00:56.32"/></SPLITS></RESULT><RESULT eventid="39" heatid="430" lane="8" points="161" resultid="3209" swimtime="00:01:34.90"><SPLITS><SPLIT distance="50" swimtime="00:00:45.94"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="583" birthdate="2012-01-01" firstname="Marie" gender="F" lastname="Grundler" license="437647"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="27" heatid="264" lane="4" points="369" resultid="1959" swimtime="00:00:37.61"><SPLITS/></RESULT><RESULT eventid="31" heatid="337" lane="8" points="271" resultid="2514" swimtime="00:01:39.04"><SPLITS><SPLIT distance="50" swimtime="00:00:47.10"/></SPLITS></RESULT><RESULT eventid="37" heatid="408" lane="6" points="316" resultid="3044" swimtime="00:03:01.06"><SPLITS><SPLIT distance="50" swimtime="00:00:41.33"/><SPLIT distance="150" swimtime="00:02:16.63"/></SPLITS></RESULT><RESULT eventid="39" heatid="437" lane="6" points="309" resultid="3263" swimtime="00:01:16.48"><SPLITS><SPLIT distance="50" swimtime="00:00:35.96"/></SPLITS></RESULT></RESULTS></ATHLETE></ATHLETES><RELAYS/></CLUB><CLUB code="7265" name="NawaRo Straubing" nation="GER" region="02" shortname="Straubin" type="CLUB"><CONTACT city="Straubing" country="GER" email="martin.mn.nickles@t-online.de" name="Nickles, Martin" phone="+499421989848" street="Pfaffenmünsterstr. 21c" zip="93415"/><OFFICIALS/><ATHLETES><ATHLETE athleteid="165" birthdate="2012-01-01" firstname="Kimberly Melissa" gender="F" lastname="Salva" license="442948"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="22" lane="2" points="423" resultid="165" swimtime="00:00:39.01"><SPLITS/></RESULT><RESULT eventid="3" heatid="48" lane="3" points="408" resultid="361" swimtime="00:05:18.59"><SPLITS><SPLIT distance="100" swimtime="00:01:14.53"/><SPLIT distance="200" swimtime="00:02:36.31"/><SPLIT distance="300" swimtime="00:03:59.34"/></SPLITS></RESULT><RESULT eventid="9" heatid="124" lane="6" points="453" resultid="941" swimtime="00:00:30.80"><SPLITS/></RESULT><RESULT eventid="17" heatid="231" lane="1" points="404" resultid="1740" swimtime="00:10:55.27"><SPLITS><SPLIT distance="100" swimtime="00:01:14.97"/><SPLIT distance="200" swimtime="00:02:37.66"/><SPLIT distance="300" swimtime="00:04:00.80"/><SPLIT distance="400" swimtime="00:05:23.92"/><SPLIT distance="500" swimtime="00:06:47.74"/><SPLIT distance="600" swimtime="00:08:12.24"/><SPLIT distance="700" swimtime="00:09:36.27"/></SPLITS></RESULT><RESULT eventid="29" heatid="302" lane="5" points="438" resultid="2249" swimtime="00:02:28.74"><SPLITS><SPLIT distance="50" swimtime="00:00:34.41"/><SPLIT distance="100" swimtime="00:01:12.67"/><SPLIT distance="150" swimtime="00:01:52.32"/></SPLITS></RESULT><RESULT eventid="39" heatid="445" lane="8" points="451" resultid="3328" swimtime="00:01:07.39"><SPLITS><SPLIT distance="50" swimtime="00:00:33.44"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="287" birthdate="2011-01-01" firstname="Szemen" gender="M" lastname="Matyuhin" license="423598"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="38" lane="5" points="410" resultid="287" swimtime="00:00:34.91"><SPLITS/></RESULT><RESULT eventid="8" heatid="100" lane="2" points="411" resultid="750" swimtime="00:02:49.35"><SPLITS><SPLIT distance="50" swimtime="00:00:37.95"/><SPLIT distance="100" swimtime="00:01:21.01"/><SPLIT distance="150" swimtime="00:02:05.64"/></SPLITS></RESULT><RESULT eventid="10" heatid="150" lane="3" points="397" resultid="1132" swimtime="00:00:28.43"><SPLITS/></RESULT><RESULT eventid="12" heatid="187" lane="7" points="386" resultid="1418" swimtime="00:02:36.44"><SPLITS><SPLIT distance="50" swimtime="00:00:33.65"/><SPLIT distance="100" swimtime="00:01:15.98"/><SPLIT distance="150" swimtime="00:02:01.14"/></SPLITS></RESULT><RESULT eventid="28" heatid="284" lane="6" points="309" resultid="2113" swimtime="00:00:35.06"><SPLITS/></RESULT><RESULT eventid="32" heatid="354" lane="4" points="452" resultid="2638" swimtime="00:01:14.09"><SPLITS><SPLIT distance="50" swimtime="00:00:34.93"/></SPLITS></RESULT><RESULT eventid="36" heatid="394" lane="6" points="332" resultid="2939" swimtime="00:00:32.16"><SPLITS/></RESULT><RESULT eventid="42" heatid="480" lane="8" points="399" resultid="3591" swimtime="00:05:31.19"><SPLITS><SPLIT distance="50" swimtime="00:00:35.34"/><SPLIT distance="100" swimtime="00:01:18.20"/><SPLIT distance="150" swimtime="00:02:02.40"/><SPLIT distance="200" swimtime="00:02:44.18"/><SPLIT distance="250" swimtime="00:03:31.82"/><SPLIT distance="300" swimtime="00:04:17.32"/><SPLIT distance="350" swimtime="00:04:56.21"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="393" birthdate="2014-01-01" firstname="Sandro Riccardo" gender="M" lastname="Salva" license="450278"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="55" lane="7" points="227" resultid="416" swimtime="00:06:00.68"><SPLITS><SPLIT distance="100" swimtime="00:01:26.28"/><SPLIT distance="200" swimtime="00:02:58.81"/><SPLIT distance="300" swimtime="00:04:31.62"/></SPLITS></RESULT><RESULT eventid="12" heatid="178" lane="6" points="206" resultid="1347" swimtime="00:03:12.95"><SPLITS><SPLIT distance="50" swimtime="00:00:42.80"/><SPLIT distance="100" swimtime="00:01:33.28"/><SPLIT distance="150" swimtime="00:02:31.74"/></SPLITS></RESULT><RESULT eventid="14" heatid="217" lane="6" points="188" resultid="1648" swimtime="00:01:29.99"><SPLITS><SPLIT distance="50" swimtime="00:00:44.25"/></SPLITS></RESULT><RESULT eventid="20" heatid="236" lane="4" resultid="1772" swimtime="00:00:59.28"><SPLITS/></RESULT><RESULT eventid="30" heatid="316" lane="4" points="221" resultid="2353" swimtime="00:02:48.64"><SPLITS><SPLIT distance="50" swimtime="00:00:38.32"/><SPLIT distance="100" swimtime="00:01:20.97"/><SPLIT distance="150" swimtime="00:02:05.75"/></SPLITS></RESULT><RESULT eventid="38" heatid="415" lane="3" points="205" resultid="3093" swimtime="00:03:09.66"><SPLITS><SPLIT distance="50" swimtime="00:00:46.71"/><SPLIT distance="100" swimtime="00:01:35.57"/><SPLIT distance="150" swimtime="00:02:24.69"/></SPLITS></RESULT><RESULT eventid="40" heatid="461" lane="1" points="233" resultid="3444" swimtime="00:01:16.15"><SPLITS><SPLIT distance="50" swimtime="00:00:37.06"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="426" birthdate="2010-01-01" firstname="Alexander" gender="M" lastname="Kaspers" license="418237"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="4" heatid="60" lane="8" points="374" resultid="455" swimtime="00:05:05.33"><SPLITS><SPLIT distance="100" swimtime="00:01:09.94"/><SPLIT distance="200" swimtime="00:02:27.05"/><SPLIT distance="300" swimtime="00:03:46.40"/></SPLITS></RESULT><RESULT eventid="10" heatid="148" lane="3" points="337" resultid="1116" swimtime="00:00:30.04"><SPLITS/></RESULT><RESULT eventid="12" heatid="185" lane="8" points="358" resultid="1403" swimtime="00:02:40.47"><SPLITS><SPLIT distance="50" swimtime="00:00:34.89"/><SPLIT distance="100" swimtime="00:01:16.36"/><SPLIT distance="150" swimtime="00:02:05.32"/></SPLITS></RESULT><RESULT eventid="16" heatid="228" lane="7" points="353" resultid="1724" swimtime="00:20:31.61"><SPLITS><SPLIT distance="100" swimtime="00:01:12.38"/><SPLIT distance="200" swimtime="00:02:33.79"/><SPLIT distance="300" swimtime="00:03:56.94"/><SPLIT distance="400" swimtime="00:05:21.38"/><SPLIT distance="500" swimtime="00:06:46.65"/><SPLIT distance="600" swimtime="00:08:11.13"/><SPLIT distance="700" swimtime="00:09:35.27"/><SPLIT distance="800" swimtime="00:10:59.08"/><SPLIT distance="900" swimtime="00:12:21.92"/><SPLIT distance="1000" swimtime="00:13:44.43"/><SPLIT distance="1100" swimtime="00:15:07.40"/><SPLIT distance="1200" swimtime="00:16:29.05"/><SPLIT distance="1300" swimtime="00:17:51.39"/><SPLIT distance="1400" swimtime="00:19:13.70"/></SPLITS></RESULT><RESULT eventid="34" heatid="361" lane="6" points="284" resultid="2687" swimtime="00:02:47.81"><SPLITS><SPLIT distance="50" swimtime="00:00:34.81"/><SPLIT distance="100" swimtime="00:01:17.34"/><SPLIT distance="150" swimtime="00:02:02.83"/></SPLITS></RESULT><RESULT eventid="36" heatid="393" lane="5" points="303" resultid="2930" swimtime="00:00:33.13"><SPLITS/></RESULT><RESULT eventid="42" heatid="479" lane="3" points="325" resultid="3580" swimtime="00:05:54.52"><SPLITS><SPLIT distance="50" swimtime="00:00:37.34"/><SPLIT distance="100" swimtime="00:01:22.93"/><SPLIT distance="150" swimtime="00:02:10.25"/><SPLIT distance="200" swimtime="00:02:55.05"/><SPLIT distance="250" swimtime="00:03:46.62"/><SPLIT distance="300" swimtime="00:04:37.59"/><SPLIT distance="350" swimtime="00:05:17.11"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="461" birthdate="2008-01-01" firstname="Johanna" gender="F" lastname="Trisl" license="390302"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="5" heatid="70" lane="7" points="444" resultid="526" swimtime="00:01:12.67"><SPLITS><SPLIT distance="50" swimtime="00:00:33.33"/></SPLITS></RESULT><RESULT eventid="13" heatid="207" lane="4" points="450" resultid="1571" swimtime="00:01:14.92"><SPLITS><SPLIT distance="50" swimtime="00:00:36.31"/></SPLITS></RESULT><RESULT eventid="27" heatid="270" lane="8" points="412" resultid="2010" swimtime="00:00:36.25"><SPLITS/></RESULT><RESULT eventid="37" heatid="410" lane="8" points="439" resultid="3062" swimtime="00:02:42.21"><SPLITS><SPLIT distance="50" swimtime="00:00:38.16"/><SPLIT distance="100" swimtime="00:01:18.11"/><SPLIT distance="150" swimtime="00:02:01.69"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="462" birthdate="2009-01-01" firstname="Sofiya" gender="F" lastname="Chassovskikh" license="485427"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="5" heatid="71" lane="2" points="509" resultid="529" swimtime="00:01:09.47"><SPLITS><SPLIT distance="50" swimtime="00:00:31.81"/></SPLITS></RESULT><RESULT eventid="9" heatid="128" lane="7" points="536" resultid="973" swimtime="00:00:29.13"><SPLITS/></RESULT><RESULT eventid="13" heatid="208" lane="6" points="479" resultid="1580" swimtime="00:01:13.42"><SPLITS><SPLIT distance="50" swimtime="00:00:35.74"/></SPLITS></RESULT><RESULT eventid="27" heatid="270" lane="4" points="493" resultid="2006" swimtime="00:00:34.14"><SPLITS/></RESULT><RESULT eventid="33" heatid="359" lane="2" points="384" resultid="2668" swimtime="00:02:47.52"><SPLITS><SPLIT distance="50" swimtime="00:00:35.57"/><SPLIT distance="100" swimtime="00:01:19.29"/><SPLIT distance="150" swimtime="00:02:04.58"/></SPLITS></RESULT><RESULT eventid="35" heatid="382" lane="4" points="585" resultid="2847" swimtime="00:00:29.21"><SPLITS/></RESULT><RESULT eventid="39" heatid="449" lane="6" points="570" resultid="3355" swimtime="00:01:02.34"><SPLITS><SPLIT distance="50" swimtime="00:00:29.92"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="465" birthdate="2007-01-01" firstname="Tiffany Vanessa" gender="F" lastname="Salva" license="331446"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="5" heatid="71" lane="5" points="543" resultid="532" swimtime="00:01:08.00"><SPLITS><SPLIT distance="50" swimtime="00:00:31.23"/></SPLITS></RESULT><RESULT eventid="9" heatid="131" lane="8" points="541" resultid="996" swimtime="00:00:29.04"><SPLITS/></RESULT><RESULT eventid="33" heatid="360" lane="4" points="364" resultid="2678" swimtime="00:02:50.55"><SPLITS><SPLIT distance="50" swimtime="00:00:33.95"/><SPLIT distance="100" swimtime="00:01:15.71"/><SPLIT distance="150" swimtime="00:02:01.98"/></SPLITS></RESULT><RESULT eventid="35" heatid="382" lane="6" points="512" resultid="2849" swimtime="00:00:30.52"><SPLITS/></RESULT><RESULT eventid="39" heatid="450" lane="2" points="566" resultid="3359" swimtime="00:01:02.48"><SPLITS><SPLIT distance="50" swimtime="00:00:29.90"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="493" birthdate="2006-01-01" firstname="Johannes" gender="M" lastname="Kaspers" license="390301"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="6" heatid="78" lane="3" points="418" resultid="584" swimtime="00:01:06.10"><SPLITS><SPLIT distance="50" swimtime="00:00:30.16"/></SPLITS></RESULT><RESULT eventid="10" heatid="155" lane="8" points="428" resultid="1175" swimtime="00:00:27.73"><SPLITS/></RESULT><RESULT eventid="12" heatid="188" lane="4" points="352" resultid="1423" swimtime="00:02:41.40"><SPLITS><SPLIT distance="50" swimtime="00:00:30.34"/><SPLIT distance="100" swimtime="00:01:13.24"/><SPLIT distance="150" swimtime="00:02:00.88"/></SPLITS></RESULT><RESULT eventid="30" heatid="325" lane="7" points="414" resultid="2424" swimtime="00:02:16.79"><SPLITS><SPLIT distance="50" swimtime="00:00:28.65"/><SPLIT distance="100" swimtime="00:01:03.33"/><SPLIT distance="150" swimtime="00:01:39.87"/></SPLITS></RESULT><RESULT eventid="36" heatid="398" lane="6" points="469" resultid="2971" swimtime="00:00:28.66"><SPLITS/></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="561" birthdate="2014-01-01" firstname="Johanna Malene" gender="F" lastname="Hecht" license="455010"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="11" heatid="165" lane="3" points="306" resultid="1245" swimtime="00:03:07.05"><SPLITS><SPLIT distance="50" swimtime="00:00:41.73"/><SPLIT distance="100" swimtime="00:01:28.32"/><SPLIT distance="150" swimtime="00:02:28.24"/></SPLITS></RESULT><RESULT eventid="13" heatid="202" lane="1" points="338" resultid="1528" swimtime="00:01:22.47"><SPLITS><SPLIT distance="50" swimtime="00:00:41.86"/></SPLITS></RESULT><RESULT eventid="19" heatid="235" lane="4" resultid="1765" swimtime="00:00:51.65"><SPLITS/></RESULT><RESULT eventid="23" heatid="243" lane="3" resultid="1809" swimtime="00:00:46.89"><SPLITS/></RESULT><RESULT eventid="29" heatid="297" lane="6" points="339" resultid="2211" swimtime="00:02:42.02"><SPLITS><SPLIT distance="50" swimtime="00:00:36.45"/><SPLIT distance="100" swimtime="00:01:18.81"/><SPLIT distance="150" swimtime="00:02:00.84"/></SPLITS></RESULT><RESULT eventid="37" heatid="406" lane="3" points="337" resultid="3025" swimtime="00:02:57.13"><SPLITS><SPLIT distance="50" swimtime="00:00:42.55"/><SPLIT distance="100" swimtime="00:01:28.84"/><SPLIT distance="150" swimtime="00:02:14.71"/></SPLITS></RESULT></RESULTS></ATHLETE></ATHLETES><RELAYS/></CLUB><CLUB code="6661" name="W98 Hannover" nation="GER" region="09" shortname="Hannover" type="CLUB"><CONTACT city="Garbsen" country="GER" email="MartinaDalig@aol.com" name="Dalig, Martina" phone="05137-907977" street="Oberer Bruchweg 30" zip="30823"/><OFFICIALS/><ATHLETES><ATHLETE athleteid="182" birthdate="1996-01-01" firstname="Anne-Kathrin" gender="F" lastname="Bucher" license="281525"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="1" heatid="24" lane="4" points="669" resultid="182" swimtime="00:00:33.50"><SPLITS/></RESULT><RESULT eventid="9" heatid="130" lane="7" points="615" resultid="988" swimtime="00:00:27.82"><SPLITS/></RESULT></RESULTS></ATHLETE></ATHLETES><RELAYS/></CLUB><CLUB code="4502" name="TSV Zirndorf" nation="GER" region="02" shortname="Zirndorf" type="CLUB"><CONTACT city="Zirndorf" email="giererjoerg@aol.com" name="Gierer, Jörg" phone="0911/6002875" street="Frauenschlägerstr. 9" zip="90513"/><OFFICIALS/><ATHLETES><ATHLETE athleteid="245" birthdate="2015-01-01" firstname="Elyas" gender="M" lastname="Rückert" license="453445"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="33" lane="1" points="183" resultid="245" swimtime="00:00:45.69"><SPLITS/></RESULT><RESULT eventid="4" heatid="54" lane="3" points="149" resultid="404" swimtime="00:06:54.35"><SPLITS><SPLIT distance="100" swimtime="00:01:35.81"/><SPLIT distance="200" swimtime="00:03:23.71"/><SPLIT distance="300" swimtime="00:05:10.03"/></SPLITS></RESULT><RESULT eventid="10" heatid="140" lane="3" points="155" resultid="1054" swimtime="00:00:38.91"><SPLITS/></RESULT><RESULT eventid="14" heatid="214" lane="6" points="137" resultid="1626" swimtime="00:01:39.93"><SPLITS><SPLIT distance="50" swimtime="00:00:49.18"/></SPLITS></RESULT><RESULT eventid="32" heatid="349" lane="6" points="177" resultid="2602" swimtime="00:01:41.22"><SPLITS><SPLIT distance="50" swimtime="00:00:48.30"/></SPLITS></RESULT><RESULT eventid="38" heatid="414" lane="7" points="146" resultid="3089" swimtime="00:03:32.29"><SPLITS><SPLIT distance="50" swimtime="00:00:51.49"/><SPLIT distance="100" swimtime="00:01:46.97"/><SPLIT distance="150" swimtime="00:02:41.15"/></SPLITS></RESULT><RESULT eventid="40" heatid="455" lane="3" points="171" resultid="3400" swimtime="00:01:24.37"><SPLITS><SPLIT distance="50" swimtime="00:00:41.31"/></SPLITS></RESULT></RESULTS></ATHLETE></ATHLETES><RELAYS/></CLUB><CLUB code="7195" name="STV Pegnitz" nation="GER" region="02" shortname="StvPegni" type="CLUB"><CONTACT country="GER" email="info@koerperrezepte.de" name="Behrend, Andreas"/><OFFICIALS/><ATHLETES><ATHLETE athleteid="294" birthdate="2006-01-01" firstname="Sascha" gender="M" lastname="Bergen" license="418244"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="2" heatid="39" lane="4" points="509" resultid="294" swimtime="00:00:32.50"><SPLITS/></RESULT><RESULT eventid="8" heatid="100" lane="5" points="472" resultid="753" swimtime="00:02:41.73"><SPLITS><SPLIT distance="50" swimtime="00:00:35.66"/><SPLIT distance="100" swimtime="00:01:18.23"/><SPLIT distance="150" swimtime="00:01:59.16"/></SPLITS></RESULT><RESULT eventid="10" heatid="154" lane="6" points="461" resultid="1166" swimtime="00:00:27.05"><SPLITS/></RESULT><RESULT eventid="32" heatid="355" lane="3" points="498" resultid="2644" swimtime="00:01:11.74"><SPLITS><SPLIT distance="50" swimtime="00:00:33.73"/></SPLITS></RESULT><RESULT eventid="40" heatid="472" lane="5" points="489" resultid="3534" swimtime="00:00:59.46"><SPLITS><SPLIT distance="50" swimtime="00:00:28.11"/></SPLITS></RESULT></RESULTS></ATHLETE></ATHLETES><RELAYS/></CLUB><CLUB code="4332" name="SSV Forchheim" nation="GER" region="02" shortname="Forchhei" type="CLUB"><CONTACT city="Forchheim" country="GER" email="karsten.schmidt@ssv-forchheim.de" name="Schmidt, Karsten" phone="09191/3512338" street="Kiefernstr. 7" zip="91301"/><OFFICIALS/><ATHLETES><ATHLETE athleteid="343" birthdate="2012-01-01" firstname="Miriam" gender="F" lastname="Pieger" license="469914"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="3" heatid="47" lane="8" points="354" resultid="359" swimtime="00:05:33.87"><SPLITS><SPLIT distance="100" swimtime="00:01:16.85"/><SPLIT distance="200" swimtime="00:02:43.60"/><SPLIT distance="300" swimtime="00:04:11.17"/></SPLITS></RESULT><RESULT eventid="9" heatid="120" lane="1" points="346" resultid="904" swimtime="00:00:33.69"><SPLITS/></RESULT><RESULT eventid="11" heatid="167" lane="6" points="361" resultid="1264" swimtime="00:02:56.97"><SPLITS><SPLIT distance="50" swimtime="00:00:38.39"/><SPLIT distance="100" swimtime="00:01:24.77"/><SPLIT distance="150" swimtime="00:02:18.50"/></SPLITS></RESULT><RESULT eventid="13" heatid="204" lane="2" points="377" resultid="1545" swimtime="00:01:19.46"><SPLITS><SPLIT distance="50" swimtime="00:00:38.07"/></SPLITS></RESULT></RESULTS></ATHLETE><ATHLETE athleteid="481" birthdate="2011-01-01" firstname="Peter" gender="M" lastname="Ujvari" license="451870"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="6" heatid="75" lane="4" resultid="562" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="12" heatid="184" lane="8" resultid="1395" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="14" heatid="221" lane="6" resultid="1679" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="28" heatid="282" lane="5" resultid="2097" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="36" heatid="392" lane="3" resultid="2920" status="DNS" swimtime="NT"><SPLITS/></RESULT><RESULT eventid="38" heatid="418" lane="7" resultid="3119" status="DNS" swimtime="NT"><SPLITS/></RESULT></RESULTS></ATHLETE></ATHLETES><RELAYS/></CLUB><CLUB code="2538" name="TSG Backnang" nation="GER" region="18" shortname="Backnang" type="CLUB"><CONTACT city="Auenwald" country="GER" email="schwimmwart-tsgbacknang@web.de" name="Meyer, Anja" phone="0173/4922745" street="Forststr. 10" zip="71549"/><OFFICIALS/><ATHLETES><ATHLETE athleteid="525" birthdate="2010-01-01" firstname="Pia" gender="F" lastname="Jelica" license="440148"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="9" heatid="123" lane="5" points="425" resultid="932" swimtime="00:00:31.47"><SPLITS/></RESULT><RESULT eventid="17" heatid="231" lane="5" points="425" resultid="1744" swimtime="00:10:44.44"><SPLITS><SPLIT distance="100" swimtime="00:01:12.95"/><SPLIT distance="200" swimtime="00:02:32.69"/><SPLIT distance="300" swimtime="00:03:54.32"/><SPLIT distance="400" swimtime="00:05:16.99"/><SPLIT distance="500" swimtime="00:06:39.41"/><SPLIT distance="600" swimtime="00:08:02.10"/><SPLIT distance="700" swimtime="00:09:24.47"/></SPLITS></RESULT></RESULTS></ATHLETE></ATHLETES><RELAYS/></CLUB><CLUB code="4298" name="SC Zwiesel" nation="GER" region="02" shortname="Zwiesel" type="CLUB"><CONTACT city="Bischofsmais" country="GER" email="kontakt@sczwieselschwimmen.de" name="Wernick, Kerstin" phone="0151/25309534" street="Ortsstr. 4" zip="94253"/><OFFICIALS/><ATHLETES><ATHLETE athleteid="569" birthdate="2008-01-01" firstname="Simon" gender="M" lastname="Süß" license="368646"><HANDICAP/><ENTRIES/><RESULTS><RESULT eventid="16" heatid="229" lane="6" points="475" resultid="1730" swimtime="00:18:35.89"><SPLITS><SPLIT distance="100" swimtime="00:01:08.98"/><SPLIT distance="200" swimtime="00:02:20.66"/><SPLIT distance="300" swimtime="00:03:33.05"/><SPLIT distance="400" swimtime="00:04:46.85"/><SPLIT distance="500" swimtime="00:06:01.14"/><SPLIT distance="600" swimtime="00:07:16.55"/><SPLIT distance="700" swimtime="00:08:31.08"/><SPLIT distance="800" swimtime="00:09:45.99"/><SPLIT distance="900" swimtime="00:11:01.14"/><SPLIT distance="1000" swimtime="00:12:16.89"/><SPLIT distance="1100" swimtime="00:13:32.65"/><SPLIT distance="1200" swimtime="00:14:49.35"/><SPLIT distance="1300" swimtime="00:16:05.71"/><SPLIT distance="1400" swimtime="00:17:21.49"/></SPLITS></RESULT></RESULTS></ATHLETE></ATHLETES><RELAYS/></CLUB></CLUBS></MEET></MEETS><TIMESTANDARDLISTS/></LENEX>
